PK   p�?X;q��  �N    cirkitFile.json՝M��F������TT�d�Ƴ{�av1�I� I�bl��e�-{��[	��[A�O�ZG��Q/&�oU�ħɾ����W�}[������ɭ�7�w�~��y���f�a{_v����û��'����ۇv�ܷ�z��c��&�����mS��b�i��r��<�&+�B�u�ܾ~{��
bV���
���V�P�f�B�3�U!ԥ������`U���`U���`U���`U�e7J�D� ���b7K�D��ۥY"R��,)�i��v�4KD
�m�%"��8���n�f����{�Y"Rؽ�,)����;3�w�%"��;����f�Ha�N�D��{�Y"Rؽ�,)��i��5��;����f�Ha�N�D� �t�w�v�4KD
�w�%"��;����f�Ha�N�D��{�Y"ԅ�;����f�Ha�N�D��{�Y"R '9��Yؽ�,)��i��v�4KD
�w�%"��;��.��i��v�4KD
�w�%"��;����f�H\"�{gi�N�D��{�Y"Rؽ�,)��i�ue�N�D��{�Y"Rؽ�'�a���O���.�.�����o�����}��QNX:��=��v�?����CL�y�I��n�u1-$4�E(��j�n�y�^��F���%l܅�;J',]�36v;�N�t�rV֫j5�-�y�^O��*L�Vf�j���2/��΍)��a�ٰ�tҧ;�UY�|�ZOW��Ӣ�b����t�g"�E�\/�����;J',]\���+�ءt����	���J',]�gl�fl�P:a�B=gc7gc��	K��;�NX:��^�õ�'0�ށ	Ǐ�i��j.k�kX>����W8~p���	̧����+�O`>���\m�|��=�p������O���W,��|z_:?��`���;������'0���Ok���'0��b���,��|���}]����\dp���	̧{^�����'0��ց��,��|���\�|��)8~p���	̧{������'0��J���,��|�����?X>��t' ?��`���=�p������Ow_��oТ�Ђ��?r��`����p������O������O`>�e��?X>��t4?��`��ӝ�p������O����+�����Ow�����O`>� ��?X>����?��`����p���V��(������O`>�w��?X>���S?��`���#p������O������O`>���Ư���O`>�H��?X>����?��`���.@p������O�����O`>�Ǐ�mNo7���?J��`���nWp������O�t����O`>�0��?X>���7�
�?X>����?��`���~tp�����+|#���6%�N�6����᧽OGצ��'5%�;�6*9�����᧭AG?��9r�i3αg�Xc��s6v�1i{�;ޘ{��y�o@��W7��Nf_�1�{���~a������w�����Lom�uO��f۶E����=Tj�x�o�� ���?��Ó���F��=�h��o�[d^b��9�-o=�sMl�j��,��\k8y���-����C����ë���Æ�4|�/���eb\[��X��n��a�M�|�/g�v��[P�xc_Xr��7��%w���i?m�1�.����Ϙ�g�~��î^��v���g��A�H�?���ͷ	%t~b� ���C	��"H(��ABA�\�
:�3D�PЕC	]!0D�P�EC	�nY$�ڜmc�-�qSJ�[�AL�wfޔR�֚�߂8��51Ąy�`&N)�n�1a>�a>N)��ƀ���7� �|<�|�R
�i}�	���qJ)t� &��3��)��]&��0�0��Bw9*�1�1���!�ĝI�N�`>�c>N)i3 �	���qJI��`L��瘏SJ�\c�|��|�R�& ���㔒6����s��Iq����)%mT�1a>^`>N)�z�	���qJI7~c�~0/1��t�2Ƅ�x��8��i1&��&wy���qJI7QbL�����SJ��c�|��|�R�Mi����CJ�7���U�U�c������wDU�/��Ca���F&��;�x��k�O�6�`\=X{7�C�z�s���i�&��������ba�zڑ�������u�K\O;�0�`ָFq��i&����Ӟ.�*WVqa�i�\���������
�ՃU\X��`�����r�Z���'�NU�S��Sw�O�%>�������>����\hŇV����O�B+>�z�Ol}�0Z��=>����\hŇV�b��֧s�Z�S�[��̅V|huo�Ol}�2Z��=>>|�2Z�սJ>����\hŇV�\���銘�%1��,��2��̅V|hu�Ol}�2Z�ս|>����\hŇV�$��֧.s�Z�[�[��̅V|hu��Ol}�2Z�ս�>����\hŇV���ܘ�S��Њ��=���O]�B+>����'�>u�����^p��:ݭ�t��O]���e�O]�B+>��7�'�>u����j�����e.��C��|b�S��Њ��|���O]�B+>�ڻ�'�>u����j��>u����j/����e.��C�=Q|b�S��Њ��v�O]�B+>�ڣ�'�N;ɜ����e�O]V��e.��C�=�|b�S��Њ��>�O]�B+>����'�>u����j/*����e.��C�=�\b[��e.��C���|b�S��Њ��8�O]�B+>�ګ�'�>u����j�9����e.��C���|b���é͇O]V��e�O]�B+>����'�>u����jOF����e.��C��%}b�S��Њ���t�m�S��Њ����O]�B+>�ڳ�'�>u����>?$�
�6�|3ݔ�bZHh��PT��rݬ�|�����s�G����2�Mv��@�*]��vaaP�=Re���H��~�#U:H�T��<6��e�w衯ce��z��X&��`:V���~?Ա2L=�s��uY<oBh+��S����XC��+��Y��Xd�,z�X&����8V������u/zzೌ�W�j>[N�f���U�6�̦�l�e^V�qUsi�NR�k9��r����_s�UY�|�ZOW��Ӣ���|9�n�L�|�^d�W{I*rͰ�T�k~��ru�LR�j3I*W]&I��$�\�)�T�ZL��U�I�:(y�:L��՟u����W{i2L__��\�'�d�$���Ks=&��zZ��N�>��Csh'���u�?F���þ�{	8��0�P���
�܅AB��"H(ts*B	�n~F� ����$�uB	�n�AB�[� D�P8����\��m̷3nJ)���݂�7���S�	�o��R
�e3Äy�`&N)�ゞa�|<�|�R
�R�a�������qJ)ϟ3L��g��SJ�xf�a�|<�|�R
�k����R8^a�q��s��)%�#�1qgR�S)��瘏SJ��	c�|<�|�R��B��9�㔒����0/0���
Ƅ�x��8���:0&�8wR���qJI�*`L����SJ��c�|��|�R�}�إ��K��)%ݧ�1a>^b>N)�X�����]��|��|�R�����%�㔒�Ø0�0��tƄ�x�������V��|��qK�*.�����>>Z����������V���*.����U�U��z��k��\��k��D��U\X�:�%��v*H<XŅ5�Q\��k��D��U\XC��B��q�`�P�z�Ъ`\=XŅ5Խ�)�*WVqa�{�}
��˅V|h��f��:U]Ne�O�%>���T^.��C�����֧�r�Z�g�'�>������>����\hŇV�0��֧s�Z݋�[�j̅V|huO�Ol}*2Z�ս1>����\hŇV���\X��\hŇV�*��֧.s�Z�s�[�+bN��|�̧.�|�2Z��=p>����\hŇV����֧.s�Zݓ�[��̅V|huo�Ol}�2Z��=�>����\hŇV����֧.s�Zݳ�sc�O]�B+>����'�>u�����j����e.��C�{�}b�t����>uY�S��>u������|����e.��C�=|b�S��Њ��J���O]�B+>����'�>u����j�
����e.��C�=8\b[��e.��C��D|b�S��Њ��D�O]�B+>����'�>u����j���:�$s�J�S�>uY�S��Њ���O]�B+>����'�>u����j'����e.��C���|b�S��Њ���r�m�S��Њ���O]�B+>����'�>u����j�6����e.��C�=�|b�S��Њ����S��6>uY�S��>u����j/C����e.��C�=}b�S��Њ����O]�B+>��#�%��O]�B+>����'�>u����j�R����e.��F����*��L��tS��i!��.BQMW�u����j�7C�a�2Лv��@7ّ*}�G�t��2�+{��@w�*��G�t��2��yl�A��d��C_��0�;�hձ2L=�t���C�	+�d���8��@�d��S*��0Y<�,ȱ2L=qq���C�5;�2Y<���gY���|����z=-V�0mZ�M��24"˼��뫚$���*I���iU�!_���U!崨��2_Χ�<�/��z�]�K��ո$�\�K�
��6��r�e�T��L��U�IR�j1I*W&-��e���j/M���뫽4&�����d����K�a���j/M�e����k�����������f�q�o�wͪ]���z�_�����ז�����i��7gQ�vSʢYN�f%�bY���z���e�Z�٬)��a)>�9q"6�@�b�h�&��#�|�1�֩�-K˧�?�S���S'.�-'�L:7����6�\L?���O��%�}��'�Q������}�~�K�\����y�ud����g�H�{�����cq����^�N����E�?bI`���Ib] �\3����e�|�%��-�+' ����k�r�K�������3���~&�K@��;X��z�K�f�~����Csh'�_���l��Vv��v=������������㟲l��#�Y"tW|�f��]12R�%Bw��Ha��+#�Y"tW��f��]13R�%Bw��Ha��;#�Y"��Ym�pO�>��@��x���x� &j��˦V�G0R�F8^��r ^*���5��ұ����S�F8^��r�QbA
�i��]#ﶴr ~�~j���=���f���5��S+��v�p���ZJ~�~j�Ю� Q�%>�9�v��p ~�~j�Ў� �9�v�$p ~Z ~j��� ��v�|
p�L��������5��$��i��]C������5�[pz���S��va8 ?-?�khw/���
E\����Ԯ�� �OK�O�ڹ� ���Ԯ�a �O+�O�㻸��qz�6+&=��z�r�N��?���kdg�#���|�{�̟�����C������ꥣ�>~��1���Ə����V�3�}�^�Uc8{=W����/.F�����?/�'0_\4����N5~^�O`�P�ڤrzH�X>��B�k���!�c��u��)��ď��Ooj���t�
M�7d�1�k�H�������PhB���!]���B�M�t�&�Po@�cHW%0�Єz�4C�2�	�&�����	L(4�޴Nǐ�P`B�	��{:�t�
M�����t�
M���u
L(4�nҠc�_O�/��uJF�)]���B��:�t�
M�{��u
L(4�nJ�cH�)0�Є����!]���B�f0:�t�
M����u
L(4�n£����PhB�@Hǐ�S`B�	u�#C�N�	�&ԍ�t���:%�딜�S`B�	u�,C�N�	�&�;t�:&�P7*�1���PhB�dMǐ�S`B�	u�8C�N�	�&���p�N�	�&ԍ�t�:&�P�
�1���PhBm�@ǐ�S`B�	��C|'
���S
�N)�:&�P�h�1���PhBm Bǐ�S`B�	�y	C�N�	�&��+t�:&�P���1,�:&�P��1���PhBm�Cǐ�S`B�	��C�N�	�&�&It�:&�P<�1�w�����:��딒�S`B�	��C�N�	�&Ԧ`t�:&�P��1���PhBm�ǰ���PhBm$Gǐ�S`B�	�	C�N�	��ȧ��"�}0�q|����F����k�U�z}PG���/9��wt��^���υ7��9�	�D�XkJ��6V����ǐ���V�p��6V���ݓ�N>���S���+,zִ�auTY��Y���Xk���4V�����$���~�2���Y���L�Irg~6Y�$w�W�����WG>j�·�4�LtL*I.K��$�c����4���$���'�R��Nv��sI�[Ғ͜��%M���7M�����ji֤��VK�0˥	X���,ͧ����<��7���u}��Q1��&)�����DW�:�[�W�R�;��f�������G�*z����G�.z�� ����:m��LGd:"����tD�#r'�Q!a2��ǁ)��}>����<������I�8"�XjPC�b:9sr��O��%N��OSXb�YV:��r�&q�i9	ԇ�L�Xu%.q�4b	Mn���ZNg��6��Nn8xa���C}�,�;���IL��=�I����^��/O/��ʧ���K��KU�%yzI�/eO/e:+5ww����l�7��n�p��'��������6�+����A�G�/��ÿ5�?u��~����m7���p��ү<~ʇ�~{�s��}�^����L~i��O�B��{��F�I���w����kԝ�n���6������}�.��/�o��q�oד�CČa|��?n���q��/�<��~����$���a{��b^O�y�jV�U��|�me��"����~�,��Og�W5�a5mB��Ηy��Y9+
�P�������ӗ�I\����Q(i%s3��Q�92N?��v��k��׈]f��ŋn�����^ȆF�������lhD54�!C/��j>0���(�F#�:y!�«p�1tI;n��W%��zy��$�4��<Mo6K����q��:p\/���%����99p\/E��e��q�>s���<�{{���q��}񦉼�_�8�Yg�lޭF��)b�l���ß~�_?��I��"���B���q���Ţx��~~�����W`y���1k�i�(�i%�jZD��ڦ��H�8�J�Ӊc��xߟ:�e�(�1E��E��fǿ�kn�1W�����a�Qm�(/V�f���2U���Kx�&Yw�\�Y�]�V�ǅY�q2뎋�V>����������J�P>X>��̟ ��y1t`yT����P�:*�W�7����C.f'_����_��q�L8��X���t�^����9��z��w�8�=��,���ϕ���K���7��Yͦ�l7�l�\N�U3����r^���M�ܤ�vi�[�/=�@7k��k����+տ^��9Z@���]�vt^�ǩ?�}W�N�����]ީD9��w���wz�l~��N#��������f��]���i���s�~���>h%��M��n�fr�f��8K������ML�f�i{��{���vj�������a'�o>�e�����a��?���uڟ޼y3ѳ
���/���1?��޾���ʍ碷�z�Gܜ;��c�V�E����<yӷ��L>ǔ�:}�MmE�O.��ؓ�p�<���7�N�X�����S�/�����z��˫�,�k�M�@�H�,��,4��oˢ�f2!$e�ׇ�g���_��RK͢v�Y�v%)�Ү��'���A76�������7��W�sH�k�?�
iU,�͆L�4�I�6gG�Ì���,)=�>�+��}�3�����u>=F-�Ӯ0����W�#P�E����S�%�ׇeC������<iW���ɿ1yF���s�vl�|}������azz���t���H<l(y�����5�v�m�t�Ş����m�k���v�<���C��<��PK   p�?X����V5 GH /   images/553717b1-fb1f-43bb-91a8-4009c3c39665.pngl{P\A����A��;�wwww�����������[�����(�^1L���=����f�~H"���  $i)1%  j  σ�����.��"�*��X�0��pR��  q����RE4��"��lo��n�d
pwwg���v66t0e�w2O��� � �ž�xd���{(�/<�5u�|u'صb�ĕc����FG��B���r�g�+q�u�11U���-l88�U�cS��z��2�+W�#
X������x�������7�<����;[��TR�n.?	�+��H ��Ve�|jL����}9̃�B�B���0��{�v���k�ч"�  k������s!���4X�2��:�����!�I���"���%�fe������2��w�����
������Љ4x� ��Rw��[��W���>�el����$�>�	Lǭ��E��p(�q��N����gm�A0`�;ʰ�G�
m%kC�20��_���c�k�D�;�\ǦCx�
���@�M���]�\ ���&#��:�ی�U�]� �L��~�Q��s���2����@��p��Ou���	�G84��8��w�
�E8�)��k�!`�n��x�$�=���P]4�5J�)%�Ԁ'�c�j�/��<������z�Ĥ13��i3��4���I� lq ��VE�5g�Y�_4^}�g���s�n;TQ��B`W�ֿɜ81G$-�C������n~�����z!Z̴��Rwl*���E�C�Q����ț>�q�!N�C�'AYx�o�+D�V�w��B�k�rq	zy!_��V ���0O?T��-��ҳ���9uj�d�
�х��Q���+�������T�lj��Q�"-��4U(�˜:.Qk$w���%��Bc����>�r���ηʟ,B�	�ؓ�����ey?�Tn'I�$��qj��S�Ggg����#-5`op]� �	��edwzϕ��ęUHhh2NNl444X8�o�>��9j���c8�؟����vv��l�����55����!cbB���<:�GF���M�Ρ���#Dbʎ��wB#"B�����p����iimUTW}{�I��P��R�����vHv&2���ۉ?�3,V, �*��p��Q$�����������s�o�b�$J:�V�Q���8�)}�������Z�$}������/�IH��
�`��-/CxS-((/�:x����qG��
�z�j��f�
+�7�:|��OAs*O*�\�Z�{��p����B! ��$\�Ł !,�ߐZX� �XֆOI�܍��*��fJ%���g��<�t�����!&�ha�ۛ��iPâ�Kna�x?G��BH�̊~�Z�7A���I{�F�>Ng"���v8���͸�&�A��in/�Ǧ�����r��?���$#�����.8�����̴�g�5Fӑ�ۭ�D�Z�6�I��\�An�� �Y�+>�ڗ������R2̎mj�� ���)0�gʛ��111�Z�6��������;��ls@�fJ���l����Si�A�<Ԅ���Ǫ�`�{��k�~��b�x�����m��V�sf� ����F��xzF~��]^*� ��O����:�25�Kg�����5��QK��#��zp" La�뛖���ҷ�k��D@JQc��e��=Q?yЅ��w�� 8����V�H�j���: R{x#�ҁ��V]i���ߐ
P�Z��)^ݸ��x��0ftj�%��(���	#� �-�]�!>��0�4i$�*�Ξ}�3I�%�@R��%�#)@5�#�z.P�J8[%a$�9G�
�NO?xwfhZ���ŪN�l�"�s��8�e9�'�������Z4v��VX-Ѽ�ݷhGU��a�W�$���]��L5��q���p�T�|x�^pq+��f�n^mpֳ��@�3�Ǧ�����X���RW�a�(q8��T	}G�v���27��s6�� �;��v�V��?���>ާN�ԆX���f��� ?vP�ӧ�+K�Q:5W�lB*j��N���F�\�c
�Wh;�"����۟�Դ�\�]�XJ�8 Q	�/ej�����Qj2�4����������]jA�	:5uE���R��e"V��ujRK��c<���ql'Y�F��'Rͧc��5���h�a���u�H}p��*�?!��ZrB4{,9o��>��8���c�V��}����KԶ:��S��Ծ>y��T� ��˺�.������)]��p��{ �������n���)�Ҥ�Äez�b3)�y�/6����y�t.��_Hg�����4p)�8`���Z��������IS�������⇢��y��^&���y��?4�.D ��	}Y,�e���i����̕��Qfff.՚�4خ��}}Xw��.��1rG D�	�VԨv��WB���?H��,�+(��K	�-��`$*�U�cL�U�jP�#�x���������\����0=0�/�;�<�;���ŞUL�n��ji�h�I*K��l�Pe-6g�a��Yx�E�pO�4;�
��v8l���G-��xȁ�1P͇��<�w*��#̋Ϭ�1�(�l�l��~�B9SugpKԳ��I	y�>d��'ׯ�y�e��H�=p��[�;�e��d\K����
��!��.���
l\�
�V�� �r����;��^J���g��%��] V��bcbc��
]<|#�����ڤMf�X�[|Xx�;n������o=���-Jӛ<$'ˮ�s�}�9�m�P�ʎ.��=�A�ro\.o+I%����B�j��\���I	���Qv_2�Skkٔ�?�)T�dЋA�g�KВ7eq�䢍_��R��R���������>�'\��}镥��w��h|��Wv��P�{� �^�Db����@ίyZ[_��HH�Ɨ��. R�	YS�*�#H�K���tSԭJ���lN{�37���ҫ���F���rv�*��o�/������Uƃ�6+u�W�i
zz����osKUn?uiHl�5���=��"`�wu���A�(��
|'�
����Ӟ��#c���c�F;��͘�l?����(̐���������t��@@k+��X��Ϭbaa����}�ڰ"�B�*M<��F1�qI���!8Ƞ��_��9��&��k����&�Ɨ�rj��(���I��No�s����dO��S��nJ8�� p���>��ʂ�҈≟�&�W���6��}s���&]N: q7�k�?_� ��Kq=R��5��+�����s�� t���K����j��5l8�X�	{^���-,��-�_`��"z)� |;4y�lhh/'%.�Pm_�ϊ�7
�^Pqty���k���Vw�W|>�&��G�%��=Q�e�x`�cC���ѩ�\����W
��s�3y��GaDZ(���"���Q4� �<C���<e�=�X�&�GNoBeOz_��
x?�mhp��~xx ��gf�����w�O�	N���?�oU6���&g`@bMEd``@�짦��%�LA��0K �����Ӷ
@¡x�m�Q�/$��yu4Tf�A;ww�������ȝ��II9ee����~�2�d�RՀ ������e 	c<W�-��7��ЬS�Q>��4���}}(��|2���R��?�G�(��;x|8*ql�q{xU�I��e��o�P)f�g`"�He�����5�9���sQBd�̓�i�D�`�KĚ*�v�E�����v_B��v'�_��Uپ�$/X�,)�7�4k	TQ�]\(��ۆ�M3��v��h���}^O�z��u.��bY���Wu0��c��BZ�{��|B��\Us�G��I�ن�m>y�JF�}��wu��>���m��yx��[
Z�L~x I�>{�?#�� -
������x't� ���e�3?1�v<�|�Ї�J�����(EM���ȈS��o
� 6�wo�V��g�@���k���;�����N$���id�^f���w}�%�2ڬ�-��c���ԭ�.�60y���xW�����ƈd�8��ۣ{/Я��U��U=�l����r-���M�@��ю�F�6�V0�d�V��A�gք��+a�k�͚6���x}��d;� wS]2X=���s�w�tՀ��"UӪui�H��AL�{	LS��[Ǜ�p�	����H�'q�.��SR�н�۹0]v\����t��b�������ړQ�j�z˩��K���;^�gP_�t�����n��&cv'8M�?�6����"�Lȭ�����)�L�_mU1j1oͼ���ē��l|�4�9�	�2�K�<[�M�̖0`0cb�֕��m�w�~��'� ���KN>��h`S{Z�N�`�e�]d�	xtW����j�y����\��2�>�#�ı"n�?� H ���p�ȏ� �.ä�OXEzC5��>n��%�y�_����}�=�3hL:80;[�G QAp��ӓ�B��F��E�m�؅6sdV6���P���޸Ə�tҚ"/[�Tʺ=�~� g���'�C����)}��`knq{VF�r["�Gp"�Т,)G�ό�ZX�I�o����%~li�h�s�ki�=YnN��M��ˊJ �g��݌"�[�D� ̙�O7��<��(�gJ���o��0����,y�UnI֖I���Z��>�˅w� ��/K�EG�KK��>�E����F���M6�c��N&��_ ��UMa�	��'d�����y����(�!ۊ8�_6M�!�]���,R�kM:|�Y�(1�ʵB��)��d�v�rDA��<�}vH���>1�`���g�	��rh{XeN��huc`Ǐb�G����-�_����E�
w��WJ�	��������4�dkee��vR��t���i/l�|��������f�����B������q,�m��o����ɠ?�i��/�v�����3G��
����CP[��x�%%��u���,.�O�?5�QKT������wզn5�ܖ��XY�>�EZ�/,��̢j[����C�rҧ�ʕ��4�!j�"�j�A}���uK�:�v�Y�t5��}�ZY ��Hidr�9h^�IS�Xj��R�3�x��h���Ƭ�%��=��C+Sx~rq\o�.��ͪޣ��:���|��3;m�XnR�}�V���������8���Q��1#�R�|�J���n^J�����y�"	�ţ�DD��Ibw���oF$t��@�ւ���E��`RW�%%zs���fT,�evDD�Dr	���q�k�r��v�D���:�:�
�˭ǃ��T��
G��!�to����Õ����i�����,�]z'�%�
5��_�
ixOO���K�Y+Z�A����<E"��h`h򸰩�l��B�1�vd|vvl\\��f��]��5�Z�Nx.Y����>��պ�it�r������|�������Ia���XO>�/'tC&� �w||,���t���z���� �"���zW�;�PPj�q������������ؠw@����W����{�o�8�d؟{V��9
 ��Ь,=���@ ̺ ���[^�f�ʋ�W]NG��ye{;�v�]�B�6:z`4���@t����T��"�v�Mw��ڭ�Hڻ��n��z��Gp��D\�+�*�7/o����H�BI���)Y�r�ƈ*Z��S��}fl����� ~zF�lDo����ȋ�߫&E{��^���Op�&]�o�v�J���ﱮ�k�_��V��[���H�|�,R	uR����������$����#�D��y��޵L�\�������F�E��I�Z�F����M��C�k�d�c��F�tXn��J�I�:��"��,�kHRA~_q���`q�D0TT���lD/X���J[9W���	�*��P6���7u��Ԋ��~�5�o���I�sb���n|%�G��G��^9C�\�P��4[h?�PQ�,!ٳ�t���)U�`���EM]RRRa�!�:��"�ٽ!��<A�t[ �T�T�����ʹ��wo�
��N�6L�r6�D�p1����v	�?s*�s���r��;�_ˑ�t��e�Q�@Z�YYטd�t��\u3V|�S����N����lP���0K��Ҧ�a�	N�.#6vp��*@�Z�"QM�F�"+�����E�� ���^���(b_	�ϑ��1޺r��B4r\4��l�n*r��'x���':g%��r���c!brwD��#�E��f��l�_���Mp����]�u�s��P=�VN�ܧ���SO� �^0;�G��N@��h0 �PD33_�afh9x��)p�/�ZhX$ \Y�Ǌ5�>�����t�[�}�Γ�+*��s��?]$M�KH����F���Ka�D��hb@��W �h��R�PR��]}5���������	yZo��Egq�&�b�tPC~�Kmuz^�b>ݾ#|8����	ž㹐A�C�r
Qf� ��x��AH�������}(���x���q��L��sG�{��� 2h����l٘�E��9}��j����"����:׿Mu��!�{��8�� a�քV����B{zoʁ��P�{��:�Fɗя@ex(]��:FG��,�m��L�s3Q����NkmaQ���WA����'Sy���y����D63)�i�T�1n�r���T�+�)
q�C�]�嬑��KIgX:�[�m�1q�{;��o�*%���u��O����q�����?�s��̧�ǎʅ}�=�x\�>��?:G=M=�mz���N�h Zq�Z���H�٩�Yq}�5Šb��#�����OD�$%�.s�}�ι|lQ�5f�D�l�%j�d��� �`���ǁ;��pf�ĸ]4��3����K�h�_��i���SĆ���lyrU��9Z�������$L�����	p7�$B�Dl>n�~w�MӜ5��P�fM�K�vj/-��
J=��m��0!A!9^ ���'C�٪��&Ey�l΄j��v�, X\N���R���q��U���D�X��l��w=�q��ƺfHF;Ǐ�G��=�͛>[Kh)-|$���xd�߀�`�oh�6��q51�h�`�$��!��jNF��_�}7��D��CIo��`k�~�_�֜"�
�}d:���Y�ZфN���ļ�գ�e�/4���)iOM�C�okH|Ǉ	!�
�r�#�^����(����z�Y�.P?�Iď�[���j+�:��$��G����9��屙c�%�=ah�
���׿�`H|P�~�,�!�ۣ�?���y~�#ԃ�l�Eg��"�NG��'#W��]�1����t�qsڔ�w4�2m��ȣ�����4d�e����;��9\k�'�f�	�E1��_�P� M�8�w�� ���.t� 10\(^�oKzQZÄL��T��\�ȴq�~o>���aaaU+K����oO�tIJr�b6r�=��x��@���i�?��_�Wy:�Syě���)��U�N[TY�R��MKz����n`�C}�۔(��/�K����?o5I�B��������%sV����c�N{k���vP�O���n�Ў$�l�\P)c���Q㧐F�)�]䬵C�{�sq:��I6<��鍦�5u�׳���\����E9��f��%!���#�n��y��--P���3�P��P�ywH�� ^"/:"
��B�-��Nv` ���rl��(P������u���M�KIש���/�J�Z��W�0�r>����JQ�6�z���E�V�늋��s+)[��{l�KkK�f$ v��K_</1�I� �����:�/N����߁�n�7��_�}��~]����m�}�)%�o�aw�B��3�K���qy'DĨ�������� ���O�6����?U���[{�IQ�cP$�7)�r@rw.HM_Q]��Ugt-�����d۾�,�~u���W�L4R�\T�C��aH��}Ƹh��=���A�l^��4�C#��B�^F��8�e�!�,#AU�罽�� �I�KsA9����y7�/&Ȁ�1=%�꡿��Њ��qmJ�����2�����ڜ���4��8���$
�	����Ke��3��-�����Wɓ6�����q�K��3��ć����1��qW�iZ_�t<9
d��26H6'�4���ؘ�P.50.�Pȏ�����'q8X��X�ύ�����X:
K���]�A����\������ݍYNI����?�RV�Bn.[��v�j�v�TU��7�3�({�����cC�6<�bk��pT���8��J0 ?�hVn�~��&H�u�đ0�	c��K�(ꙣ $���ŀ��B��������~�I�Pu}_ש9Zp0��_�ݯE;��lhlV�������v�hG!�׊)��m��9�g���l���������5�����ݚ:rRPR�qp`I�~�����gQD�G1h�l�a3���F�6D�����./d�D�����BY��ª�a��F@"���� ����>�B˳���#l�������TS�law��B1�娉�c�Ȼ���+��f
2�R]�0�V(�&�`�콴f���9�!��+�~�I�k��RPO��4ח���}C��3�Uf�l�*����]�cl�����ҩ��=�����>��� �l~��E`Z�������G��'�<p��1O�BUS<�`j8cy���h300m�!��ޣT���vG\����̯�1�ԑJ�̴o�Uum�bMu�8��Ǎ��tt�
��8wf�Fx�O���V,���i��璁���$��IM�8ч�:�V�-��o&�z����lP�Z�?o����E�����d�B��@k����:�=>Yh�Ϊ��ڢ�l�o��(��"�0
�C�"�6ReW]��a��YZ�*J�	~w2cݻ8����y���Et~C����X0�(x����8��4`��"z�
���PH�M�CN���U�=��vʮ���Н�	��X�汼�U��7�']���9�af�$Ix�MA��Ҟ�#�P�%m����"�\\(�4-1��"B���n�$�MY���/��sX/  777�=]�[90	��	O��o�'/yE� [Zm����zF�u�C�r����s�T�C!�u��Z6�<����B��~le_$�ϗ��ꝰ�4\��*睾ѓn�`��/r��l�#�p&�1s������l�K�F�@���g���g������f�
}x��	b��QWLR�s��0V�E�����}���]	.�XK�/s>:��\t�)�`ؿ�s�>yX������@}46����l�PF���\��(�.O>����k��o;ŽT���_�
'���8oy�?<������B���L��K���nU%3�=�Is����}Z��B�\f����â�鸸�%�:jZ���ҿ�T�����L�/��܄ϖABy�H��c�� j�c���+�������;�m���<Zo�7x��2����ۋN���`%Eo6\@t*�����bf����;94��������:��})�#ޖ4����	h1�CG�(�L9I:�'2"�E���_SYَ�v�'�U�z��Y��eGOWk�����/��EMMMuI|����X���h�۠�KZ�41���
��u������:H>�� �GS����(ɹ��G���l:�]�#��
&Am�5C����Z�h�����Л���ľҎj���7Xd2�GGj�H�DI�F&�
�=%���T�P����ӧ�Mo2��$�M��(����ߩ�Rx=1_wN
�F�ij.֌�	�oV1y*3��X8)!~����5	�O�o5+�&e!�x�x���r��v8�����ZS#�"���۬�ç2����}���z��L���|c���b����xH�>���IH�sZ�Ľ��
�
� O���� Y��m�OO3������Xz����f��3Ƈ.������^�i�myy�s3�Q�D�
)�4r�m�:E����r���zKW}���wO_	'���r�7.��������z��M��&l�	�������E1~�;<8j'�G$�x'��jqe�CB�
�Q�5𴄺�g%��lx�9&k��)�(����"�%c)n�'3�#���8�pM{�@���7\vT6��tB/���Ek��������;����C��Xw{����
1�*(H�2�ڗ�mؕ�ԣb��nv����F鋒³Q�J����Z�N�<�\D՚WƟ�7�מI�gu�?B�N��i�pu��K����_]_��q6�OS$����qF���fP��P�JK@��`6���d��:��$&f��]?����!��n�n���L�R������� H�4���*��QU"n,��G�B�ڞo��X�����%�����EwS.����!����3���sݮ�S**86�I�B��gK�[�F*�nTH!���nmcs)�v��|��\)��'K�)��/�Wtq�I�5�n������`˭���ڗ�Qᚚ_�+k|��& �S�(=�c��L�����5�C�]o�w�z\��,�����y��/��{��Ξ����(��V�Vrӵ��a@�G�M�J;W��Z��.ټ�lk�J��~��Srs�h��T�A5��h���K�������j���$1qL��>  G�LS�����k��bG���>��h`R�PZ��ԣ{�%^vz�԰R�*@���RI���{0��Z�:�f\��ʋV^��Ǎ�k4X��E��J�i��wZv�N��=�jdʌ{����$K�߸�yuu6I�y�+��G�*N���1C,�_0ыvZ��j��4eyö�O����(�e�I�\r%m����x���D8x����֏���w���bڞ��;��-�`��$t��܇��i�H])}�x[��2Z�!C���}Yd�������撥��sXB����ٲ�KZ_�
j��XY�D�(�Si������Ru��k������(r|�R�=����E%b��WBs�}��G�;�������j�vc�l%/^D%KՄ��RF�y+9X��eB�A��᳧��1�]�-�E�9Iˇ~#-�<8�U���ɔ  �	IO�Ҳ<�CJ�Oҽ�QS#oֹ����WߔwMʗz��A��:��0�� #%R�L��q���u�f%��_W�Ob{�Ij�ɦ�A�����"~ ϔʮ��dcu��r��	磡�=����yv�/���c���q�w�PS�u��JJ���]M��n>���E4{}�0��d�!!�9�8±��G[��Q�!g02���j���WᙜT���/l���K��x�|�=؋"����BAA!\D��#��z�����0Tϊ=ԡ�0�� ���2��jfq��rQ}1٬�(Kv���'� 5���|��������`��+>�Y�������>��'a�E��U��w��6@0�h���eg���ݵ��^��f�\���UȜ/��{������n�$����y�*<�������˝�T��5�����y�&�2���?����«���w���rM�%p2����bY/�Ç�ࡃhEܬ&�j�ݿ����:*��흂���}'\�,�u�>#�(29�x}���s�C���ţc�/�ɣ�P�*d"*��Za�g����{s��e�;9W3�i��~��¶���p44�2���L�M���l��ҡ�7im���j�n��Y����Ǒ��4��Piv��$e9Lݯ�W���vr~�M5�Է݄f��Ԋ�E32F��_.�%Y���r.^�`�[��߬>2��W'�����2�rm;D���%�ms�Q�_���u&��E�3Y��l�&�8�o�p��+���v�� ��Ѳ�2n<�.����(��c4�R3jN�%A�O�]���nώ?{(R�g��|tEa��9bd&����Z���-Ώx���<΂�F,�K-*�"&M�H.:�8 ��_���l���mU�a�@?}.���vt	�$_�2���t��\��ZRv=��VĤGKY�L��F�[���x)�����#��O"S��c����	c�+���а����� �S�k� �!0z�s �pL��~xǠb�{��ѭ��e1쁴��h�t�����N7Zm��J�^�P�r4$���b|�K��0kɎ��v����|8����y8��ߓ��6��A���98�w�(�H��;c�}�f��~l]d��hId�sYZ�+��(�R�3���!�|-��d�A|��{����-�y��>�N�%������޸�ek+�������� �� qR����HL��h
z�-9ͪ�NZ⒐�֪Zj�o���o��,�{���"\�Gm8��r�-��~/�U�Z_~��0u��mŚ������� ������"+� R�M��TQi,3^"W>�*oH��g:�\A��Е�Đ%X�4�oS�gt��)3����d�F���W��⾓V�^t���wk<N����]JGmd����M����������F������ˎ�*�Lӈ����%�Q�㦓s�ܖBס)��2{߲Z`�]��Se� �}��'�ĩ¸!_B�*խ($�C2{��0&ov��Z5ܺ�j�����(�f;swe��^�&�HQaR"�26�v�j�S7���L�i�^���x�딡�A.MR_�O��C����''���W��V`%a�+;9!`.dr֟;q�zK
[r�sw�|-�EN��5�_�7kz�F�+B�*�\MB�|&�4��������S��^�����v�~E
�J��b���9�e%}Q���&��Ҷ��î�L�t����<֟9�e#W�ݑvo���*@@T���7�sτ����/D�X��B$#d-\˲^?~hst���V'T�7�g �}7_�G��ѱg��� ��P3�-m*�8��s1+�vxq�5t�߻X��;�TR�Z��w%^�tO
�ܜ�ſ��+ec�3--A�l���<^wJ���H�2���VVVv�<�((�nn�j�z�KK_�ng�otOd�u�^;��p�-��/�jpH�+��4ѳ����\|��26��Vju��V\��2�,���A	�_@@���*nD� qW�:��������ֹ��D����!yǷ�:���I������>�W�LL������7�6��fޕ4��v;����ÓH�D�9R�,T�eL���v��H����K�M�Fl'�5����Ҧ�t�j�!�M�E�O�񖪊�C'���o_)�_(����&� GJ}?��~:Hq�B�c�� R�*��K�9�K��O�T�D��U?h�xLk&9�v��F��Nn��Υ䟇������0WW[1�FA=�����`�	e�aLnCE�ktl#L�����
s#���oA��Ԃ����/%fL���--π�»��Wi�H59m�.:�E\[畘����'h�`�Rg��L%A����y�u��`g�D�� �*��˝����s��JJ"u�q!TWW��Y=D���1B�FD>2�`�ab��x�����B"X�<�t���j�m
���
����M�66��Q��$�}5��~~Ё�
�����-)��o|��6��٣������:>�����⟇PV��C����"l�$6K�iϰ�} ?숦�׉.>�~[�"�ߧ-I�_W_ϊD�e����證���w_�m��<�W<Jx��N�Fܹ2��y�Y�� )�����\�ޗO ��'�,	Ou3ۣ�;_$f33g��	w�ZD��]��A����uw�U�<l�Ə�j<Z_qyfh����#���Ak^��ַ�i!���m�EsI�V���%!�U��7:�d�k���^��`>�'������/��]H�~�/��Ǩ��	��h����8!��D�u�_������F������or9F�|�?�l�rw\\if��c-�/>�B�r÷�B${5���@��X�d�s;�*����{�AP��St��`��w�@<At��!6�۠��s��{�2��ֹYg����ME)f8N��ǡx�BÈ�a��xmWW�O�����TJF�T�Q�g:R��	�Ζ~��S��_�u��k���L�`�����A�i-w��� 7��R�Gs�7�a�9Q�3�qև�Y�r����{+�ՕV�WU�*�6�3��Ë�<6ฃһ4}&�>��`�Э\�����XǑ��=e\��֙wz}�V��P�G����=\5�R�R�1ق+r�FBӕ?��օ��?���y��D�_\ai6G�3@�.�߄�'Е�6������K�0�=
���d�Y]JA{��X �u��������+8�x/7��H69ȺfO��ե7��@-ϴݟ=�5
|��n6�	�����]CW�i�՚�婺R}"����:#��?��**�M��+G����C �Ƭ�&E��պ<ޥP��6�R���#Mg����iT��ZY�.`-I�Ϳ<�+C��w��A9��JY:�߷sMP�͟����kuC��rff�de���n�m;���e��1��q6��8�P*��V�2UtѴ\S��)p�k�f
�e��7�R�/��󫄣�a`o]� 1d>m�r������*�g����-`��:�q	۠a��q�-��+�ۜ�{?���`����(���*��xz(��v/6�krqw��{zzj=�-�� �
�������r��txThBrD��!D~��#�M���+�trs}��:q�t�� AP�
j{�D�{Ƚ���; ��Ω�ɟ��sq�gbvP�[][[���G�;2�]�δ�Hp8y��f7Et�ڲj8��.FE7#x��~pv6��k�8���Uڛ�Tlg�{�^Ht|<�����?
�g,MO����
�T��j#�F^�:8�眲�-�K����ݯkԈ.l�`�_�Nx�MMM�g��E7�!����2��8̻�m�	��ԩ<��F��0���G��T��ط}��h ���[��c�@�{��N�`W�(0��,+x��*@�lx�*�j�M߀6?S�����m�峤x����ݛk�\��9Y���D�9�w��O��딉QT�z�dddd|BB`C�Or2r��J����o��|�z�!3ׯ�6��n�eI��� ��H��[ B2�Б�K(�Zh"��ܑ�3���S'P��ȸ��a���A>nbM�-ߕ��j�h:��]��m��FHX��O��"g�ˬ�>3�U�hʌ��-��|��G'5ɔ3uh k��%߹��(�zʂ-���Ή�̈?��BΌm�5�Z ��\�P/���b?�
@5��C�ϱ-�
 �� -��-m��kP�ܳ�R�;k�?�Č뗺�M�U�T��+3��B���\ݬ9[6�~Ⲿ�hf�98V��3G���;f־l�����A�7�޻�����H��Udgw�$�V�G�4y��0y'3�O���|��ٹ�f��l��D��ԓ$�'$
q���Be��{Cuj�m��ny��UjO\����X���Wd�4I|"����'��bˠ��K���(�8����w�2��j���$h�P+: 2 �8�Q���������H� V����-��5���X�G�Z��EaM:Ȋ�Uv�tF�O:E:A����6��`f�3wyMA�M�+����t�
�O5~�O�l��<UK�-kV����#6��<5���;��)��1|�s���L��ӵi�f��������õ��Qc"�	^����e�m_��4=ok۲��k�<�^ c`Q��py^v^�0������cc.˪?�2��y��{���#��ׂv6	���b��B9Ģ��U/��v�N�W��-5&�~V�M�����S|;%����l!��T1�����w�2C@KSHp�Bybߛ�$����1����t��b4��a+-�����⪱�7��	�bR�X��EE�Ӳ�N3Oڝ-՜5e��X�*�^��B2^/"�Z���1���h�5ƢtJ��*�;r�(�#��F�`��~�bI.B��, �r���X�J���EE�i�d �w�ǂ��f��)g��p7_n�����߸:��1�?�@'���!&�8���vS�h�۞����n~�p��'B5��
zݑF����?�������0��N�^aX/���_�C�k%����:~<��%L3&�������$ғ��:���ׇ�����~��Dw1�9���\�&O�_��o�mj/�H�֗f�I��l^|i�v�s:M�X��
YK`��Z!�7���;��6l	>9,U�O�&�R	��-�y}9�7�x�E�^�|hϚj�S>�������C����� *;�C���8�f	���zV�(B�����n�5�<�G��H�xa�P��{bT�b����YXP������X���������i�q�ܰ��M�V-�hA�6�H
�cWb����j���lТ��g��w��qk��}�fX��]�� �<;PjP]��j�������T���N�~�z��b���h��!G�+�\ĳ���|�6#�|QH�u���#��ܧ#(��2�~��\�I��v[���@q�Tg�"pz�����UʴV(:�6���V���z3V�C �f.�	݂����o��k��I�����iؤ�ڸqҰqc�Nc��m5�m۶�o��>����̬����`���ꬸ��X�L
�mzq�ԗ��}\�#�ϟ�iQ��~��^7�wEb�H��a��|=#i�A�p'���?Ek�|��� �oZ��@���Bg�7�A���fP�P�����ۯ��$7�	ڞx\\\�)�8�b����Ju�S�U5Ե��_��y"��scy޶[Awm/W�6N&��Z����K[��x������o���x��_��"#�.����:���'��y�������M�Q&U�|�����73��_0�3�)@�,�Y�Jf�jD]��Y�B�)
�d��Gw�-?���]t�&-߇��	k��ENx�������Y���Q���J��ױ�L���yJB%�� �������38��a�3bqd�Mu~�tv�l��j�p\����D֚*)�~T��#�]�6?�7[`sE�u�*=�Đ_�����9�R�-�*�z��Y����be@�K���2��<��y����a�Aw$w�u��Sp��X�A����׼N��B��M�
�\K�� LL�_ ����o��ɉd/��uR���@%�G���F�:���fFmo5���z
<��V ��U���=�"�Kzq*#Vzzܰx���i�o���:P@���ᓍik��G&:f�Ka�7Q9sx����1D�z�Uu��A�̢�jb]]������/  �a5���b��c����'�.~rQB@��r�z���_�.���z�����R������f�~kw��ˬ��B?�asS`���k��o���ӧ��|�j⓵�D�o�&oI\�� !��S3mʓu�C]�T���˞��>[cf6�k�0&Y��L�+5��	$dk:���ԜϘ�c�eLDI&��PƧ�(��4Y��tGf�m�+����y�kH�&0��pvK�l�l��ԍ��v��r�2Cs�a�����"b���լՏ����N}��χ�W��ݕ�=.�/U����ڠ������n��}3*l��y�k�U|޴��Gb�K�s�(�����3���gV���8�z��}_R���'�l��v���U���,�.�����ܱ%�4C���2�ק�t 򃦸�x;+5`�d˓�$���Ԙ6��c�<��;x]�fm#�=�>ܷ��>�3�j�5*ox\�����B�b�L��l����%�	U�0�뼟�Dh�-]l�l���d��:k�ksW�]㎲6�W�1@�K� ��h�����sѝR2"�	�{w��@9O�ˊ2�=/�fTO����/�����p!I4FaԄ��܏'����d�����y� m��.2�~%��uʉu�&s�-	��I�qT�=��\���ҊL�������KǶ�a��#ƛA�e?����B�q(��+�@�x]ݯ���-0��C��2��\�j�b���mئ�b�-I;����#��"��o1ZȺ!� �Za���.���;��DJ:Tc��FP���k�-	'[�~��?��=F���w�}��\���v�\�_��J'��;Ñ����Wr.�Xy��G�ߣ�hg$S��e�ax?�K,|��J�(�x@��]%<`
ܞ5��r.���hy�N;=��vϧ��P��Hi2;�t�m.�g�����q�hN��۾��f���g9�m �<�>�3��D������57?�{�����2�{�)jrr�jy��J_Y�1���0��l_����y��a���ŭâ�YK��������*��No��ٲtV+�L��kNe���<ҥ�~.�5�&�ؗ��F�Yk ��5�&$�B4��%:�~�T�s�O�*��re44[��֙�#�>8�y�e��1��r��� ��1W�`�Aֽ��ih�� x޲��H�Y���@
qĐ{Xq�H��7ϓ0����_~x�c�ܨ������5>@;{�eG}�eO�b5�ݺl����1\�� �r.P���`�/�(�kuL���[����Zt��w����rv�Tkzhi�:i#�A�sv�씠�4�PQ��ɩ�������F�uǹ��&��js����ؾO�!'u�����mΖ�"���ޞ����x�+���#ۿ~$\p����{f1����fVR6ǽdZ[�;_?;�z������'��p��g:ԏ��t��;F���ǻ��_5���6��]s�{��oph�2��
���7a��%D�\��?���}i����Hm����x�03g��q�<��8�<�y��J1�/G�1�ٕcJ�^��������(�!fa�"%��l����T����wC���KT���v��{�Ȑ��K�R��F�d�x|Me���dz���w�.mťŤ�U{��fo����CC�Qk�|MRT,umm�[qN�ʊ��l|���N<��zO���vA7<�:%}קOP�ā�a-��*����56WAq;�{b"�������v�Rt�SQ�l���.y��[��T� ~zfb�a#�-h+9��Z�^P�@커Ƹ��_��2�H�:WR���7) _v��6�><ߟ5�1P!�/����E�(��&[Kr��&}����F*�[}�2��gcs�!��^q���ysv6a�U�)�i2����њ�Q	���o���X�?/��|���N7��?��l�Ean�:����E�RrfL�OVt1�1���=��2�qRc�R��Irc�L�R���b*h���p	��Y��h�M��Ƕ������S�T�Ӧ��N)���NP}�l�R���_��^��

ak^���?ۍ��u��G��G�:��h~�p�����\e�ܦ����ȸ�҂��S&A����e��|�h�S��ނ��&zv���Tb�8��`�ǭ�j*�ϬSȗK�#�C��u��5^E��Qi�~��y[��҇��\:���A�*mk���(
�� ��v���R�Dd��)6Ts�|r�O����m� ċ{����|Z���܇'���NA��:cs���'ȏ���?i�+�3<�o����&�m��?%3�?�!��9�bA�8�^�g��Tv���L�N�D=�7'$��p��:�Ĭ�#''����)P#҅/�h�D�S�ū�m��6�ӱ5C�]������?�����$�#��;����,l�����	�
��L�*|�rY�r���K����=�x�}m5������V�2� --����B�d�Tƻq�]a�J���Ctu{[i�U���č��P�,�����W�FH���a�D�)!����
q˩MY]͆�r�Ӽ����������^�;k|C�sY"g��D�P�u��y��x"7x���1�����l����t�#!I~�L=���Oi��/�ރ���.��v{ �]�������G�N+�9���tr4�.,�y�{��H'�+���K�����Zy?��=�"��Z�5�?���������<q�d��mxU_LD�pm�rk_M��Mο"[O��
w��u"�殁��:3���ځ�v�5i�S���2V�G
JS�]+��cfXu��愙�_hu���K'%�VW�X)�������s|6wg�G�����J1�Բ��(�6��a2T�;�S�������rk��g���'Ɲd�ZX�ё��u�Q�~�IP7�传\�����q�`�&/�9˳����#��zz��`3Ե�Lo9����+�f��_B�u�%��OPQQ�hFz�,��X)����i^�\�*��۷\=?�_|�NL�;YR?<�U�kҝ̖����ofd&q���@��N��%�H�	���'5��˛kV�-��l�{�@�^U�C�l�ѝ�L���'
*�Ё�"d�b-Z�ٕ�-��B��z��t�J�둌�����_WGG���;ӑd�\���%3v��C�B�_��Y2R���|Mr%135�|͗��|]��B5I���'������t������h<�0�z111���mfi)"ۿ��Ϙ�~5'b��ДC�Ԥ��Ē��DW�M���μ��%�U��@ti�J�����|u������D9�x�d���%�mk+i�2��� �8>R�C���_��f����nX)���*!�S�/�͕���w�G�q�(�`�ќ���
��6�oWE�_�����T0��"�=� l��'���t`�+�����N��g쉙@D��M^�(H���w���6��s9�_���p5��P|����EDjhBU�ba�1886v�)��1��B�v2�����s�w��N�I�����XTa��ĩ��?�:3;35��ݿ�14��*�|YM��������I�V�Q˅�x�{wNHL�Q�gn/1�U�I-���u)x�ѿ�h	���n7m� 9P6I��eg�Nx�p�n����5�4+aK��c����s��W:���>?/a�2���jow�I�}�L��Q<(��Į�Kֶ��Xׂ�
����lo��GPҴ���0��î��6D�S��4�o���"���8�0ԯ�ͦjo7��?�5N&@�i����$ۅ�7�=mC��T� )e��#�j]I^w6�25�isib�����5��4����ѓ)+ȁ�F��������y� MM�3��2�淕�J��&���)����AQ���Q�/�M�\��{�Պ~%:�J"'��GItP� �ܒ�aD�`�әz�W�}�TE������f����ծ��êtf �7"M"��ե	�+��1G�/�rf"xCee��g��L�R;u&���k|ڐ�l,OEE����嫙˥��C������̊���Y�μ?y�6'���~�]�kk�����Vhg�?t�[s����׬^�)N�
��Qe݅E�S���ʛ)2� 1~]]�ub@S�����4'Šu��5-��o�P>9��r4vaB���$Qw�!�w�`�	�D�|��r������]ܞaͯNke�q?G�	f�0#2D�S�h���2��W'>=W�e}uU�~�������#�o���C>w��,:M�?D�_�dR@Sr|���/Q�F�q?�bD�fs���������O���(��d�0�z!�MPo�����.�E�^烙�s#(���2#�P8Ի�$��+�'����GW؆Nrdұ=���x���J:'�
.��#�ߟ&5� m1�,x\p��$�9I��o#�������t����m�Lt.39�+���Zo��?N�x9�<���`��
��<wZb����R���6.�5��d:�e��9?����fipY��A�Y���#�]|[D\� ��7ff.:�%�0�'$��G�"��|�|��Jՙ�id]�,��8�6�����a�gv�F����"��-�ґ��f�Q�+�t�%v<k���$�ʉ��&�v}�o襥�X��%��d�ׂɡ���xmk(4���/+�Ε�^����ˡ!��
���u�&�mT��@�w�˛'+WI�<<v�c"B91II;��5Մ��4��כL��KG_���e��������3i���F�`�A��hڷ�iX�l8���������<3��+���y�!����|tOt���9]9�S� ΅dOC�����!uB�з'����T�v�»�6pI�N����i��$o^+�z3��T�����f:&>��GV�kXWV���"�}Z�ު�p���oM)�0���g7n�!�R��.�jv�ӽ�,J���!��"�\�:s�[��+%�v��L��>Z�-Rai�O$Φ���4��%Ք1��.q�)�oʐȷ̧�맪���{�R�CWz�
ֻW�"� 4�TsL�9�����[1���7�o���)���D�rtxٜ�%�(���z=�E���c��"_خ�#c�4B����D)ݣ�\���tNӿ�.$��Ԑn�o���4�~�݉	E��In�v���6-�j�#���KK�
����
r�1���|*���Y2�����B��-��� �."�ے�I�SNYI���m%�������1jZ������m��z���w���0$�!{7ԸB�`L��Z�F$���>��q���ts�Rz�����~<���,�7����zB<�҇<�Ѿ�X�@)��
���5��ۋ�����9��q��#�^�Tq�����?2E/rσ�e��V FzG� ٝ�4��� �;�a$,7�@4� ��'WC��{�%��ru���i�8�@������ 𷨊�ܜ���2�,3�Q��Nr��|�7g�o9h
��ؽ�~ߺ��u�_��(Ak)����P����!^V��:5��yAT1'���&&&�rj}8LZa��Ծ�%F�ڲ�\�+-SC;��($mɊ|�_�c}��\�^i�*b��������Z��#"H�R�|m��Y����	�۵����3s��L�h���yyLn9X�]����EGE�����U>"���Ha�Os�|G�urڂ�F�K�Rt�(�7���3�I�k�̖���ŝ���0�͜����s�Ū2Ds���F���_����I��xs�p��h�4����oM�Bv�HnY�g�,�^f�d#U����gtW�rh�K��@���:�Q0�S,W��l%�g̛�_mB�:Tj���F55JW�٫̥���B�����td��Ib���\��y�s����z�Ũam�c�[#r�`���_Ψ|&���0��Q0AN;�)�%w1���I�	U� ����o���YX\�H1�"��xdj��۰/u��|��ܿ��Ĵ���p*��#P0K�0ANr�5@�χ.. ��/���I�g�3�##���c�%���:T�R.]T3c�ͪ�bb�bc	�������3�W�^��[Ӳr�s}"q�-����S�I#hh+Tq�]&]�i�7D� T����H=�NM�0��X�����%o]Q���TM*�x%��-�I-�l$��ަ�H���Tohh�����Mb��?��m�݆�c��.�f)#c9�X���Τ�9C��P��͍ا��/���I��w9���ޱ��C$G���Ώ�;~�.�������P>�ɋq���D�׽ѡ����p'�:[��u�yV�U�74�f�Y[���ۓ@<]p3d+�-��C�t\�Z
��%�j��t�G���%M~P1�����P���SKI�j�lw`��̘�`�TXxfvv[I��8ue��-w6gkYu!��l�R�r�xd�3����cvb�ik���p۵iQ x�:XW��*�L�To��3��d6�[�����N(�P�n:Sm12�~�2*>������V=���,&��33�e�R4*��3"��`2���t,,·t��E� ���������#�����p�o�P�������ggg�'"�����%�,6���<���zj/���0[)��o�(�����r]]ae��/cP��R2<�.=�^���D)�m%����%�9\V�� !&9= 'k�m�� W��á���O����x�~�Y����C(/�.),�c�Ú��"��m�f�ƴ�U���.��V�I�wm϶l�	�%5D�|b�xa4��H�:����®�]�3�(�Té4������;de�$� Д���m͖�	�z�[�}
����Ӟ����"[j�����с�ךĀD*��$^�N�L�h2�*4�-x�8�?��P��SQ��K/��5)���T	��ތ5��eS�Z���� �����Q��VJwQɮ����&�t~����k�!��)}�ar)i��שȬ2y2 �^�ie,�T�[��Xu��.���P�_횂g�hM��lE- ����/����%nKM�򢂒<�O�6J d���ߌ@&���`���>l���(ܫ*155k�%켕��5�N�a�=M�0~�!��G��/���hMW��'����ո��iR�Ww<[��.1�{h{BP)�@{�Αg��C5��܇��d� ��n�=J��t��F8�9C��u&�臐o@rr���xQ�̲��?�9�_�VﵕFŰPPP	.ư際�۹>W�ω�o�ֆ�683��:1;19�;��k���Ғ���h���BL�*]��[:_Xi�ഽ��#`��#0�����9}=9����B��%��5��T�l�F�ʶ��۲nnk� 7�8#D� )yP��.ڙH��e&�;�[��QvN�U���{ȋ(�w��C�Ep�R�x�-�M��qf)�vZ#n�@����vw���#ڋ�m\~�F��Q+�����3&ymn�JQp������x~Ѡ�����f����Y�($ߧB��1����6SOf��٪�{T�b���#z�vLO~F�8ؠ�ٗ�)�W���"� �t�e����ɾ-/?\��U���=<,.�b�m�xC"�a@��vrr�(������:��iV��?�ol\Z����&��Ge�wπ���"��p�d�<@�bU]N.J���i��=����ۀB�N[w�6bM��7*�L��s\��ʺ��aOh7ÞMk뗆�k����R"���WZ1IJA^NZ��O�S|!�}����9ЇI�N��3�����['���Jj��u���Ĳ��b|��׿��a'�?��,���=Y
�2jD7�Wt���td�)?���=��4��Ņ�{Zg�$��]��W�S`/Su������v��}���E��m�C���ݏVw�]�05�	�`Ɂ��n�,�������H��5��ݒP��1��_�8��'
�,Y
�JEq+TF�L��݌uR����º��#-�mQD�Y��	sW�C�E���<�$�:iZ�Y����Tĝ���i��
r���x�	y���F0��ik7�U�!�	�ޟ!qpp��''%%ua���?ř�re��7�A���@��?�\��c����h�TO��h�]�w6�A1����%h~�k^F"u������v����>�P���U���b����}Nw�V�=�g2�����
�U� r���0e��,G�� �Y����kD1�U�Z��+*<��#������I���	����Fɣs�Wt7�u�P�Y:���]��(���������-��"ā�f@�?��}S�x�𧋜���/������E8�$ܬ�*�&�,+˧��^P�$Oy���mI8�g�?s����)y��B?��j~����K�>�{+%�"?C��Y�
SY ;�/�A���矋k�S�ϟ���)?O'n�����AU�#�I@e0E=s:>����d"q]�hk6=����(<B	�ab�o*��HPإ�����yIk��pTr<l�e�Η�S�OF��c���񳔣�L�5a��v !�Ƕ��N;ft#�b��Z����%%z����ۗ6W~j�~;;� Z��TxS9�H��g*�r�)�Ӕ�b��՜y�#��L	0b������9;8D��ɪ�#��)�m賨�%sSɀ�-��c�J���JLL�BXjz���y	U���gڱh�1�#59�&�c�T;:&��X�X���.AHy�PR"�҅䘒/y#l�N�n�}�N�p�����4�Z���J`��~vS�����O�r���A�o�L��G�>��^9����!;�4zH�%�|@x����|}����.����(�� 6�FE� 8|l�� ��po�_Z�g�0���VX)��n]���C��97�XĢ��kʍ�{��s|�Hm��%���XOF,'��������G�9����kl�X��E����ݮ����)nb7$a#M���wpaD���}�0e��;ڢ���֎����^h�&�Ϋ�2��夬�Ɖ�g�m#q���= �%[��C��0R q�)���)��-��1�2�6��p�i�U(��j^�ҋ��]�vp�7���W�4�C$i+M�EjM�e�^�p8?�#�����N�w��h��C w������x(�jD�ק�i��O�)*l�4�j�h��;yn;q;οO{?g�cN�F�.�Q�[<w��NVn8�;G�H�%�'�.��S��nc%6D�E�#�"B��k�IV����\�Q�v^__WYova�1��_����88�&��:����D�Zn��^��-����L�5O4�{§�����>��t��G���?i
;A>��a�����W�~�^.90� �������	Փ��jY�9��x���O��i��jN����7|dㇵ��ɬ05E���ն��۞�m���
�=2�����70R���J3cNf���k���#5a^�)e�X���U%��*��M��>��ܓaT:�`bѝ�(�W.�DJȅT Yi��a�V�ݐ+����Ͷ�1L���򽦈8����̜��>��ݝ���˚����Ռ���g
(�<Sr�}���0�$'d��3VՇJ��V�: Z�Mt��kqM�Kݞ���핥O^��OӲ?ϳ�u���t���U�NookR���qp��Z\�|1NV��3i}�Ɨ�;�N$�����+�����[����3�J�U�^�].�.W�m׵��Ǧ���g�,��b��q�2;�w&�?�?�_4�@oF��L�H�ь���6>+h���R��HǊ�ŮLe��e�ڧ�������`�m����8���m�	c�U��U�����?'2��C{��vؽ���{�p��b��sA�Ƿ
�.����B�oMUڭ����`����C?�D�O�ge�KĘ�cQ��}������.��n���x�U�ʦc��\��1�y�G�"�}����+�3�u��̂\_�	=���S2�n�1�-�E���^?8���9�� ��ꠡ-��"�h�#�W���p��P:�xZT%���$B^^�Ĝe����i����!m8^P���C���;�������wӸ<J�b|n~էWFE�V9Nk�tf�w�����s9n���$�XXX�~����Itε�_r�;���E�:hs{��u����{����
���[��,��:�dk8���7<�yR���UAh�C�&R�fpG�kj����R�d�)� $9t��!�$�{o�ާ'q�3��m�hBE����ɂzjHצG�@��^�c�]��7A�ݺ�ߗ�5%sd�o�}�~ȿ�?@A� ��yZ~�-�i��Sb�2P��@1:�$ /Ͼ|e����v�
�{r���y�Y�L:�{{�"Ķ��Ҿ�N��y�� ��"�|��i% �'����n�B���"�~� @��]L����c��f��k깸45�_6Ɔ��M8ԙ��~�ׯI���ϖ�X���&��|��h O�5�w%�I�wHUĆ
ȋj
u�/�z�U�KWqq����d{W��QaΥI���OT�=��E�pI<�^���,�-Ʊzzچ52�!;�.��jHI!����&o��]\�B�&jJѮw����3���@��Z����S�=����$6���Z/>@�_�j���T.`>�4� $gI��u�l~`m���\/̜r��)�Y��\]IF��&T��NM^��Dѻ4�K,���;1>�B���M#/w�U��_K@s	Ê��1��шTā�1���%��8���P8��\(�&s�_� ts*��2#��ZJ,�/�������q�3�����1����ژ�#T���x�����15yzr�74���Ę��6@)�4-��/]* �"HD�<�J�	Aɞ��z�[������x�_���(��;�)��C���ߤd��h��k;x��'�R��q�l����O/CC�;{	JG�v_d��X�v+����3���8��̜��k������>cv��!���[;T�A�H���3�cZE��ܸ�?s)++�~5D����ص�NN�.��iP�
�@.��oo��:,Q*Q�Y�Z(E�B���䄋�O���3_�-&���ƻ�T]�K�{(��
B;o��P��ֹ�g؁��Āi�8=E�����/HO/����r1�RgmW��/���ȃ�a/ߝB
J#rrm˶�N 3�����c�W.��T��m�w�r����H!��XT~#Q	a\��� ��qa���c�j8��WS�q�LZ������׋y��\F&��G��:���I{��p��r!�_x��������kp��/;t�rc|�jpD��ťJ�W�C����\��>���^7�>ʊ��������eύ$%�y`l&�� ���!1�P�)9��3��i0�B�Ʊm�86m[3sY�!P�l�%}����ظ�M�l��~��>�Y���	#��]��?qs�sss?���_��0�[����]���Lp�|�b���rK��4���Z_'q�;A# ܽ~��C��Q�����z��P8��#���&W4�u����i��MIM�ww�$���H%%�b���%����;����Ơ�5�Ȱ��y�g�g���^��2踈܈H�������2������*��z���.��-�)�sW�����˻/���B"*-�do�d���|�[�^���� ^�}$髼�;��t "��ߣ���������ô��)�ڞ����rK�h�=O���XJl�z�ll:�PS*W]P�/,���2 n��s�hWs�Y�%��w���V�͡յRj2""�^��6Ի7�AR���*Ftf&uNvM�����6vvfv ���Ĵ��$�'~����i�Tџ�'��6��t[֍Vyd^����=�e�B��0wg��4��t�wJ::�"��$�K�ۿY�6AYsj4XC\^^N�΂��*����^h���<��6����J�A�T��y������VVad��&�>��}KJ���T�M;��X��~ ���oo�|7[�//�*Kv���U�����0���ט�J*$++�r�O�9i�pZ���2�؃�z���Zk���F�yHl�J ��b$~mϺ=Ah��  ���xt1?gwF���hA���ŏB��0�̆#����:�O�_��z�p*cm�4�v��M)�����
��H d~ ��9�[��p�[hm��S�[@��G�65?��2�㇄�7q������6� ��W�R����F���[��eb�=C��84���8�z�����_~C��q� ��tH}s4���h�M�"�COv������IOO~��!`$�񮁡��uqu��}�n/�HR�}�LZ��r��J��q�sb�#<���F�A+8����+�����7vwg�Y��t�n� �ֆ8O|�Fy�_�*���;^��AFF~ �߾y�Y �1���+�R�vb �ԒiG�h��F:�FS��D�^?qr��Y���&~5���hv�T� �t��>|�\���ox��>��@@Gp�y�����W�VARˤvt�@UO���č�����̗9}81?/f`������c��091�2��*�%ס�"��@n3����A�|2~�Z�)X�L��iv�t`k�G��V,�W��� ��tV���� ��è��<��.\C��%�v�s��|��iW��G�)�Q�H����W�TJ���C�Ĥ��@|=��?}���hf��:�� #Uq1�u�.�����&�!�X�WX�64L�:��v�d|��:� y#~w�rr�V��������z����h24hö�A�?y����"��-l%121��͕v��6O��s�LBUUU�Wi'���T��ȯ9Az�elhCG'��x�\�^���.�Q ���.A�t�s�}q:�@���ޞ�?����8�"�
�R�_�*C�����Xm�qI�1���p|1H��)�����b��0��G`�M^��p�����ब���4��e���F�}݋����Z���H�z�M�l��Dl�664lT��wOd	m��!/�3����묷ypz�8�����C�SA����}�?����c����y �Dn�������<�P�";Ln-[��nt���~�D �����n>'XY]�2��A��&��j���~��O���v�
9q�����-OJJ*,6]Z�Y	�\�@iE{.��~�b���>���P �z"�g.���Sұ��)���ۦh===\��A  Յ1=_oU��􌍃^��}Es6�+����=�!����l�hJ^�

FG�	��X��k� r����]]�������>>>���*Բ�=���U ���$5x<����|5"���E�<���c��J���"�xrs)�<���U�����yh�r�0�e�G�ۛ���";�zC����?�&��3Ȃ�
 �s�����&M"/���g(Tz��k������������G�
a��}��3�$����v�t���F1߅6P4���\Y"�S��B��?4��˸����uM@�, A�M��	�;G_G�ʏpp��"����jq盝���׈����y|���D#Xrr2�0 �̺D�p}�l���	������c�H�������J���� F��XO� �P 2�m�7���-��n!�`��i�{�F%ZDĖ�ͨ���Cqm|u�AR*·��rr��4���.ӰU77�Uۄ����|��8q s;�n���y��M�Z�}��|�����z��l���۩������,JQQ�j�)��mOū��\8h"eb���	7�).5�̂���1K5�����AHLqqq���:Vn>�A���~pt�5[��Z�-���o��?Q���&#�|u}�e���ge���� 2V�y{}�kdt�Dvv��
�ONN2sr|� ��n#� ��3Ǯ���d����Y�ٌ���]Ê⇣�
#�y��V����:|='Q��S�����*�u�ܼ���}}}���p���߀��D"�9٧�' �i!!!A�_�~-��q��(-�?8>�Ex�'#����,���<G�B���F�h?�h�6�@X&6��|��))aKKF�e6�&s��:�!�j�ʵZC�Z]k]�֫��BO��Ɂq�Gijj����r���Bg�ݫ]���NJJ�\Z��� 4J	� Ձ��qoR��]�� D���NM��Ó~c�j ��<l�=��2��iv���T�@�(-�B���`��Ô��6���L��;}a�)��y��h ���F��--�#�l��D14�����a�������8�-���$2Ci}�`�r�4臌L@��uVJ�@9���M������rƱ����=������!)�J�Fg�P���J���ـ���ϟ?�E��&�onNA�Й��@D+�<����*(����tsc#� ��5�����Am�|����4{?'7w��*��d�Ab����f�?ț��Lg ����̂���~��=��W�]}��� ��7ce�;�Z��� �ȠY�|y�I�k��/S���Xf��=��K%p�֏^ߡ;t�Tz�����U:���Bz���:���1�?u+�]۴>��e�����f�SW�>�����
���#A��������N۝� �XY1����A+�,�P�٦�=~��Se###=mk/s+��\ISq�lf]<�!������KYsg�S8��  ����������	#�������"�i�����$S� K\B_��Q'� �v���zg������tZ�OR�}��I������
; 1��O1���ds0A�{
�+(��dЍ�M`󏈈=�ⱕn��=���
Ӱ�C)�Z˾[o�|����_�5�\o'�������Jߧ����,x��2�*`�+@ $�@�K����"\
P>P��S���Q^/��ڡHuPBJ�Р��
���hap�^?$�Q�%�_��R��e��"�|�t���Y�_�"~��6E��a��ݲUPD��#�M@���Q����h4O��8�c�eu$}5�SV������s>y��f��ëz���7y��d-���[�`�ml1��W�s���Թ�%�z�����*�Y�����؎��D�. �u�T���3�� ���Ay啘i�@pڜ���
�c�����n���e�l�X��\�dee%~��KQX�5���*|j��i+�)��vj���w~���M\6SL �m�V� ���: �Bq�� �.��SɼJ�W��g*�ԏ��j�H�"�,)���^W�����lɆ5��s�G������Q���掁���a�v� ���Y"qwP�&d�0t`�	[V"M�J���h*Wu0�hUMM�� >>M��ͅ<古�� 3�F=�.fA�曒�v�!׍��[7!�����[�����M���N�?�i6��7kR�6��A�T#���&����ӽ�=3ihj.�V˫����}�]*L��/�]0�H�'�
�Z���\mr8Xm���c7��ζ5��`���'�b0���
��_c�'42 Y�!�7� ��D���}TF2��3��3`}��Q�b����M���/ =� �
�J
U���?��"2(�#.>~@Z�h	
	�B������Eav����i�i�,f��0�νu�g$m�W���k�JUz@)���94g=�w��v��8�֦8���7m\ �[�^�J@���:.�+k_��8��T���"����+����M�.^ ۝RU�_�1��%�o �V�؛����-ѩ�o r�o��������`��~U��	`d,"��-��J�'4���[,��խL��F���E�B��i2bBBP2�p N���t$ *Èx��#�ȹk�z������
�1@�J�h?u��N���a}ӵ��b`V6J�[�(��}�H���n��dĀ4'x�	}co��3ȥdC�w+�[
ff4666��鉉J��B(��$��fgg���c�
 upq}k�N���8��10(ӧ�Ɛp�cY�����Sf9�#��H�)�ը&D,`z8ȉ�^0��H���z�*��k��-�HH��4"�tKJ�tHI���� ��)Hw7�����y������V�p��k�5��k�����}�H��:@�Օ�`�W�fgg�>O�T�� ��1[eնv��ya��[3��������!�_�{�W�E������S�'(��WR� S�<u���p�e@Y����1�}�ω�L	�jzzĨ��⋁�^�'����^#��*����{b����bx�3���s����>-bzZ�!���/���"���J�Pd0-��m����aO"�ߧk?����Ag/	}�R�6h�*:�	�}i�P�,+�ҹ���D _�JK9D���ggi��	j얈��c���,6���zU;�۠�nL���p��[���Yh��s�MÖ�|�&se`��텘�½� �+ȼ�IJ�$=8?o���ڛ0;���O��.!Whњڋ�=�HH|�q��4�ORX��U��Z.+�D��_ܯOrFS�''�¹"���JJI�pr����	� ��AH��2K�
z�?����b�Bn.Zh}v~~hG0���F����|]6 q�8��f�ی���߿_ �V��!7*���%@���!��z^$�U�H�m�12�Z����yi�̷�����]����˄�kEQ��4��/R9������##�W����$d�����L�[��ru���ʪZn���<t�1ib�Ƹ�O>B2''��P���ʔڱZ���ӭ0^��t����K(�]�������/e�F{G k*u(sp���3o"##��^�~�e��u{�ggn�
��aC��p����2��d^� P�J���7� �+^�<�(�<���I�7X��<2l	��� ZMd?5_���&u�o����~�Ҷ�z�� ��i��\�!�6�_���:!��� �U�|U�e���̤����̷�]�'�; �v�p�b������� ��2�򝀏�UJ�q�%�'lK��������z�֒B�����ut٠b�1#��Q����']��`�����@����ӎ���AFA	_|�=l���5CUg"&G.	�UfB fHx�����WUU��_��K �o� Hf�	�|�����d(


J���.?W�`����ҒLX�+�_��ߩ��S�љ{�k?56���sa���,F���;�@���e�g*a~�����R�����>�"V�.�%q�WO����/6.�A�*""�# ��0'���� J���# {���v��gVV �_|!F`ZQ �N�{@�d�4H�$:����%�xG�&�j�i>JcR���W��)܄Yc��:-��>$��5Y��(���MJ�*�o4��J�:�� ������t�N�'K�ؐB�K���*������ �?�tv���I�-���7.cN���uB��(3��V�0B/���N��X0�魧�=x B���q���8۟���`�C����R?E��շ����������>V���d��v�����_M����e�a��]�p ,!�צ��o4�/��J�'&##�|���e6���2g@� ��H屟��7��[�q�nk{}&X��,-  J�q�a�+
�]���-C�TJ��h�O�'&���P`������C��?"F��FE�)�k��W���m����1�Z����1xw�28^�i_�I�|���ɨ_�w�J�,Ǚ^���v����������jy��f;#H_�_~����!�/-z� ����X+��ڪ���hi�z��GZ�&�&�v�������7�P�\�W�������dU��I2n�	���%:nR2e�o���j��'�ڛ��2�D���=2M���M��ļ��~u���N�G@ƄQ�_�p�X"`�>�:�;�� IB f}c�y�A���;?�\p�?M RJ��i���}�u��<���"����
��3�/�쬭1���k��W�|?���q����_���3���7�����dNr�����TLF�����r��|�����S%=�'����/e-%����<v ��Yzd`x�>1z�	����$hXT|Avjj�/uEE���%�ʹ6 ` ��)_�{�.k��/l/��<��6 a8dda "
���������������4�!~@�� ���x�/m]a����-���KС:�%���wvh���G�j_n��=��{�kD�$"�ku���Vc���-#�5��r��RT��&� ����̋&�bX��i��o$�`3�EB���)�!8	������Sޭ䞴#ޓ��:��JmY5�ϝ��۷/.��٭�f(�T��׎�/��TUUC(my���|/}N���!���e��c�?�������btTrjr>�Γ�?����@�)�8�?^�BDA�O�D_6�N8 �+�9rY�v���� ���W�^�;j#V��D'���$�.�) ����y�	�0086�3i/L�am�l�8�vDD� ¼y����O�����g�5TY_?pTb|'�󬁿@c�ޛj���Td��ӹt����t��R28d+�e!J���A:�}D&f�v(4 ���,;��Yͨ ����{��3;���� Ú�@j�jW8��a�������E)�M�Pp]]]�F�+��n������k6o2�t ��d/saWJ�X	��I�}귄E6���	3�t����.h'oa#8FJFF`Q�q�W_����𻃣�=��V�����>��?Y��`�;-����ٶ��7��M�7t	��qiiQj���\F��
)������S(i�k�k6Q�b��\�h@��;B0�����L������Q��-��a20V��]����؇��M[U���0h>��o��l[Xx
 �0�WIV�2f��1tY�߀����ק������T�W��;L�vs0�ͨ\;����P*���ךz��g�o�]���ϵ|�%��=�-kkk}��jf1�%˖�̆(a��R�c��]ك0I�Ŗ/� �<Ӯ}Ľ�q���O #(��lhj�c ˠ�1�KS��5#)�����Hb���*�cP	�~#;3Z\1@���z8�DPHɟ�����E�p��b��%2$oOOO���z��D�L%x�����4~e^�SV��8�4a��]�4��Жm:����Ʊ�an��C����J��R029��~2�T�1Sa�-j��}	dvؗ���� z��FwG|}��<�	̕o�Y�NJ�G�Ӓ���s&��PFgKGC<:뷎��4�Z䵺�P�H�0J8?��I&�|h}���k\���(e����p/�ܖ m�̒
o�:]Y_�:�6��`�Tۨt4��`2O�f`���6�&эeW!��WPN��C��`�Щz��
�5V�[|��c�\��!$Y����u��;���!.u ����o9(��L@��1	��QO!�a`7_K�?��	���Ob�^��R��fH*�v�++��Ý��lU���=������6�㐳lg���ZF�m����}A�����ۃ����ͽx�t����Q|<=��nJ�;�_���U��i���H�E� ���p,m���:�q���G)���M#g�}��������η�\}��-/�p)�Q��4���B"ۦ� ���9)T�@�Ʒ��pB�ǡE��&�#���sZ�'�D]����һ�ų�V��V�KS��:Uj�ֈT	�p��p?�y�"���Q̊�����L����5q����(t�c�kjj$���III�&&� `�UWR�3�2�i��*�~�0� �s'����D@ȱʿ���fPN�r�`;_��s�(�؂��D�����~���c
8m�2l������N�����B��)o)�,kLd &��k�`V��,6�wE�YO���|�w�:���E�*�/n�`�<Y�ٵ+Q�4h�x'���P�_���#�YY��dܨ��T�_i$ ãZ����r<Y�ZH�P���`�r��R3ٯ���w|
��_�D��ө\�g�E&''��ޕ�z�ﰎ���4R�lŪS��r��}���d��T�T^^�=YLe��l��2C���,V���}nN'��%+�|geTT��xp6\<<ڊҟ?遝��'�h���vc����#�����|$��TtPv��Qm�0{r9U�i�ŔN52?Raoȷ �I�X�{��+�^��e�h*���˗J���nB#2�4�u��o<�,-х��3���=�o��5T�%we��s��o�y#��R�>�=����uhU� �˕$��*����bc�Χ��<�v�@Mh���QEJ�+**����q��=/���jQQh$�DS��T��+Y,�.wG�kV��>+������@������W=A��Sɇ�"K++rk3N�:������M�Dd�0���/N)�������KI�.*���'����w�n�RWW��K>�� :�(�c{$����z ���%�hJa� �L��7��K@�@!�ˈ������΋f�tk���QڒkU��Ĥmj��v���u�L� ���a��jXZl��Ţ+5�^}�8\��
'���~4?>x��b"C}�3���g&] �E���)Ҫ��8�!����� �(�H�ٟ�@�8(0	�`�z�(�	e�ѭw���� R*� \��j�p�L�����'���y�K�ep�7��Ćn�DhEn�Ӷ|�J�w�9����0Z`آw��X�
�#������4�q�-��YBB����h�撜=��X����f�\��9��:�G0?@�����i�<��Np���c{GG���N��J��^�җWUI��T����-E��1�����F�*� ��Q��3�^�w���w(0�B��x_�ڒ�p�W�q��E;��J���]:?]����H]�����^�.S���npp�+��^d�����Lq� �n[
?I�n�i1
\�I��}8�X-'���h�N�D��囐����"(x]]]ta�bb(|�*������[|��Z$�W�/�����:Zm�^�W��L���y�2��Z����nE��L�l����O����4e�v��42�����;Rn,}ww:��硑����7)�*@��ֱ��o�t�M�l��4	��X�*-�ZW�a0��%��s72*�E����<�h�\��&
6
���ǆ<����ߗTЅQ e�����PmB{����Ĩ���*F_�c#�������@yf�[���R��1Kg�z�wB�V2�x�Icc#tT����۰�$��������G��@L!�J��eJ�Ϸo�����O���%%}��^��о���2E���@yI�K�y�.R|b�P.��c~~>t�8�^#���#��$�O�R(e�m���7�"�;m��|�X�O��ð�̟���`�TD���Ąf�9��TAF�[[[�0�����Tw����dX����wu��#Yy{����XX<�M@W`��4b ����0�R�g����l����wc���8k>Nȧ�~�2tpWHW�xJ3լ��[��p��e-s/�}�_͋܊5�E��������JGGW^h03~:8P+���3��}�&<!0��}o?�c�<0��}<|�aD��F5##������y&
؉d�dO��qO?�Cs���L	<F�3?���

�њ::�'�}W`Ԓ]��W:�{��D-�DLdde��
� s��B�#���Fjj� ��,O���M@P�*�����_deg��$��U��<�9XS��+!����.������m��ʧX���<C���[J�^��ߒ���>�D�W"��8���s����pF���&M��xn�U��r1߿���7��O Ôh~����78\l� ZVV6^ Q�I����n@��������ʇ`'9q��M�P��|^�Lb����(iȟ�jRf3co`��E-ţ�&%$�<��Vd����+�ɋ
�����]�UR)UVm�Dv�9�H�$�D�&����y�α�6��oQiV9^����f��<t�� �d��AP�9�Fx��6��m �$k�҄1@����I���������g69^��&�� Q��|��KDcF��|v���Ӱ��tgX@霯�vK��s5���MLh��P��$���FᎴ*L3�bl9�qjh�8�y�|�|}bªרYGM�;����H����h7�@`jjk���S�������,40�nB2����RI0+������@^��`�ݵ�y؄���U7�z"�\��J [@�CE��g���u�MPk��.V��1|"O���"���7Y�����s�茶���@��𼬗g�<�����7���mUPsa��,����Ӊ��A"c��e���>��@�M���:�NE;%��Ab�Ss~�BK���;YY�΃B}��:.4� �����V?��
V�Q���I���-f�z�����Y��u�K%(S�'pQ�|��LP��}�����m���=�n�`�4 ?һ�M���A�K9qܔ���/�0:ɿǇ����[|���~(G@i��_�i�>;sZ̫���;�,m�Fmİ�s^�nIa��ڿ�;h��$�y�l�6�k�?sY��e��]?��W���x+�r��u ϫ�as�B+B�0��rb�q.5chDE�1�--6��x�P�e���=?����-�CB��t�=��;;ˎ���^RaS1�l�Ժ��46
}�g�q$�˞x�b�,��,��T;�ꐝKg��TK-��'Ж;�Mʰ��f�Rf&��)		��Ȼ?]���������7��YT���{˒��rxff����}z�YȂ��C�&�5�0��8�������2P؇ ł?�D���ǆZ��%��G�i�h��a�^j~
㴞愖�o/�ǎz�5@����u���t�Ki)GD$y.���Sg��w(4����Da�^� �H��*��ڕoK�3�{F��ۿ-&S�uysP_D�\"յa�Y�R{�N]�h�̞����I�ηD�����6�r�i=��ÉW���K`�����Ή��9��q�j�X-ޚ�=�v���=�����u�H_]1.(�ϝ�y�G�\���Q�):!�!�I�$`�R�ZLtc�qr����/������V�cb1̤�s��v>��P��<F�0��������}G\�8�)��YuxD��O�=48�@�J�]N�G!8��:g鳴�,�[�3�s�7���b���D�Kv���h��k=���7���kٖ� h�r?��Vן>}
��#��h�Zp,O ��%� I__�|V8*�����:0{񝓋�/5�) �@�&�<6R<�/ (6'!��'2�`��<�2pZ���z13��;#�g�U",?i�w����R�`��`$n��4�̲NKcf�@�>??'	�/���������������TQ���@�;q�p�~� �tz��=GY.�RF@@(����#X�ːLjmd���5���-��NĆ'�VD�� �c��s������V;Z�D�#����� � E7��_|Z9 ��[|Z��c�5J�	�r���2�v�-�"�I�����C�F�χ`�'�p���E�0�(��:G��j(Y��>Z	���o1Qɇ�;�%��\�����Q�.�1GEm�i b���[��&vǶ6.��N��)�5�Z�s��7-e�,2S����H�N����7a���nh�o�����NPG3�s����pw��\v�B�VSO�pڤ��D�N�O���hY	@����wj%ɹ���� ��>�]���������J��W��By��H���0�<F4q�B��g��B�� G��΅σA���x���qf>�ۤ�x	���hH�������G��	sv�G�g����e����l4����묹~�yyy�G��ڒv���6�4���$&��I�rp`�}������@HI�Λ)�=+���@��O&�O�E� #�*�z �'�p!�c
��ց��Wb��M��;z?1�2��-��J�9�3�����L�ul�M�Ϲcba��z�1������{�x?�]nBiۼ�v?����u��b���X*K###5[�22Ĭ�5:#cc\

L���1�����3fR5�&���~�O{���*mF��yX����d��Д���b��Y��{���{F���ў�<[�XT������{W9�\e�v���F�������2M��'��$k�M�^�l�DfQ���`��Z�=�	x��@��T�Ř�Ȏ���^�b��?�X�t���1}����||��m����=���^y�Tng� Nzt��·�XM�rA�|�^�e핃��׹~���L �Cʼ��3z���ܒ`��;��@ 
m4�����/��ta� �ʁ�	쾴\���@�y3����L�?0����m ��̕:Hj���5[���G�������W��5vx���=���_sVY�Z妖�Auϥ��~yu��|XQ��n�9ꔝ��2U N���ޞ����-L�����·����A�{Q::��>��IL�%������kݑ���/�n�de&�O-�a;"��l��L�?�0������%����7>��@�uUO@�9��dQ/j�xFt���1�P��d=T�����U��HQW�G���#����O_A���xM�_����.K�1^�L;�sE@�-�� ���Hb�	7{�)���Y	3�:�����q+j��\�@IW7i:jj��b���.�)l�'� P����+�x-�=�xE-{<	�@g8�r33��[C�(0�g�x4�rى�uŀ0Q��bbaI�l][[#����r�Kth����4��ta;�ȣ.b}J+ �����"�_�Ke�����l�0���$��-�r�xt�K��π�t��'a��vD���:-�K����ם��P������0b�i k�횯7M��^E��<�4#~,�Z�]:�j1lٿ��A��Uɕ7���3� U��x􆠠P�����o/L�:�}�]U�H���� ��}�x&66���@LB/U�����N65Wi7m����OKK���KS�o�l4��鈺���[uu�0�}�S�%��!�G
���,��T��F�u����J��ʗ<�@I��6�>����b?:Tz�h��Ʉƾ������ծpTTT�H�3 ���y'��L��)}���E��NK�|cRRXNu��b�NÊ@^_,@�(���4*�89q����?c[ɭ�#P��V�Ee6��i�nʻ2�)�i�J���SȭI:5s4�N��a�V���6U���L�]T�?	c��=��kv?ݔ�;��u
�z)�W�W�~��{5���Ӥ����ч%��"�{��Y�=���HL1'�@u(�.��E�߽{R��N��)2�JXtO���8��G���@�-..�v�* �MWYCZz�CUU���qT�FzzD}�{��O˭p�C���D��n��M#�������l��!�<��&""��7�W��j���JB���KH�7ee��q��9��I˼K+�H�w��Ӌ��*�u./�Ԅ���KJJ̿���M-��nj�psyM'R��|,-:�җ��N<�G����8+[[�7��p��|�!�'F�F4��CXA3�P�'888�z����ʪ�|J�^OPt%$��Mw�*�o1/�Ǘ]C�-�!�x�.�u<�������g��w1;�Q��1��N3����k\񑕽��@F@O�b�Qqs�o���m0eb�i�p44L��K+�����Q*S�R��g����'vpQWGh)<�[��Q�a�H�{�����ݹ�U�8a!i�u�d�7%�����Lsla��v����0�����o�猬p�7��;ܜ������H�*&��L�3��x�h�ޯ����|H�8�;1|�� G@&�b[�=����}�5�1q>..����&�Hc[5!��AO���c7L�Y�N�hTЋ�RM����V��yo�N�����}�0V���7}W�)���rj5B��/]-@����+J�r���sW<����60S$�G3ed&/��c*���QD����3N�w��?�i/�dd^��mʄ*�P� w�L�23�?ޝbC;��?L���6���g��	��t�$����+dhAS�ۀw\ll�i�p3 )�c��p�`�c|_P�ʢU�!->��ǖ�(��Sub�eǑ"_&��0s�"pב���t����C
|������ZЪ�ହnݍ1c��]O�r���Y��hy%��p��g�B��ðs��*�K���������E�|
l*>[�xu�*�	�z T��MhT�2��u�;���N��}���
��x���cZd`h����h��n�ͥ�^L!��y�#C}E�Q*���$�jE���ON��z�R)��G>��hI�S�qNۍ��1�=�J����;:�O�*��l��������_����*p��.8�]K7ɮ����R7�p�[H�^��d��Y@ms鍻�?9�K��ϱ;{�٧����7�C=�ey♾�F��/^��<��4I\U8&L���$$h�k�����!�]\\��r��|G�g����
���f��);ɳ�VS%��.�wI�:����N˵��,F\`f��]vqY�0���:����uؐU��A���3n��l�~$>oZh|��=V��%������ĮR��5|R��oK�(�m�+;;a s: }ј�����.EXxx���$"���9_/ZX��omѽ|�����0�uvv�������|J�20(�[�e'�Q���赆��(��cu�٧��-�)Zb5N.ޯ�C�����z�}�ͅk�����9̠L�㴈?3��5iϮ�&�$J���zQ��f�K�-{{�`C�GsQ37ׯ�b®lp&B�7�lkm�}�����R2�r��I�vtj���j��u��ŝ��gW��/�_UU6"��h��vS|_�HH�a�{tg�=�D:ڃہ��A$��k\�5�J�8��zT����fR�}u=Aӓ�����F����q�w���.+Kf�-�kj�/}��E(q~�qM����۾Fz��N�r�giN��g)&�{�w~F�"rr,#��,�\���푞
Z2�J-�zC/��<y���[TV��}�vK"G��T�<<U�<v��<~��8[YM]�U�c��՛��0��V�����6��ӏ�q��}y�i���6W�;��k�Ə�b�̯��x ~��I�X]]w������Y0�g��ѓh'�, ���v��r�&���MA��vc}�p�B���}�)yq�Y��"�Ă�<����yu��V��1ǵ����vy�M����A�Crx�t���pD��f��M��s�����0��<�a�6E�4v߿]]1�K�kݚ���۲��~��_��B+���ey���,���K�[���[qY�Ϫ��=ǉ�	�IG�����������9���qg�����o�&NZ�/X�h��*;8��_� �n��om�6'�}���R��Oj�&t"s�vq�S��c������
<����>y˲�0�d7l�>o]a��cz.�g9	��t���ݯs�y��L�}����%��\aW�~��6�|)((�6�^���厶��5:mvzǜ�y������	܎�y�����r�̼>C�Sg�����	������@5	r�T�����������4(�Ê�Z>;����M���A�'�"MZ�\\\$����٘�O&9_�P�
�
L�w��'ܸ+?��Hh<����,����S����<`1�gM�܆�2�\�[�|{�͹%����e=�,�|f�C!8̑n��� �������Մ����p��Ή�9#Sc�K\j�E�^_�D�&��-����>\60���V��3{YY�#.����]�/Y}SJ7VŁ��c�~�X^#�ya�m��W�2���J*��0F�/�h�C�Q=�±;��q��!��s����23Ԁ��ݟm���(.���F���W{�[���]p=[g;�*���qnvb��}�����5� �q�+cRSj5���&�*~g���+V����ݑ�x��(h�ܯ���m�@��l�"�P�$�z��BA�.���:����G�1�p#������YG�4�M̑�k{Z�uʏ��Ì��G�o�N�Ϗm#��k�}:���t�����fާ.��qdy�sݢ�����\���ԙ�!�;�ֵ��� �NM���G�l����l�pT��է�y��B�2�ܳ/�l��p�?V"O�)�ꅈ)D�]挎2��'��~b�2�O*�O����o�p��	��V�@�ſk��s�ju݈S�)y:էC�D�K��T9�J�����_��&DP�We+�����e����U�(� 뀏��5��@�B
�9%��5�\�>}�Bd��T.0�]���_V@�"Z�d�w`�߾0�G~�З���:{"�߿�|1c�7����!A��$e���W>q����9i���I��N >k��K�N�ɜ��-�������7in�^��1�{�<�����a�&��j.U��um��0=/(}�9=�(���B׺6͍,��F���ʚS����~�*�ߝ������a��/0����4"�B�j9຃�??���N�k�1��<�|X���~���T��x\���l�0G��f�o�'Ჰw��b<%K?_�#��]BY����~��|q)���&#��!�����j�g��m?����0`j�g�y�x��`�f\�OM�����ŏ�bD���{�)!�ǆ�~�kma,l6�O!�@�,�t��a�3W�Zr~S��4�@VD�c[GN+J��_���;�5��%��Ƴ}�l�/]��(�>`���_�3/�u���z��ƪȕ۹�n�	�ﰑRWA��;!�k�_
���|F��3.��,��/e~(M8��;���V��
׸'���qK�r3�Ognr{F�C�Z��`QX؛�{=���E���bflԄA��0��i5cQ��څ��K�A���^��\������UUUd���#WX�o#�<�o�J��;�)0�1��+���
����W�����*zn$.dRH��
	͚���AW�֘O(������c)������W34��=~b��2������c71����>}��oN nmő�D��篋�`��Ez"bVn0�����7�=�4�^RҷOΒP���)������'�����c�q\�QcAH���d��h�K�n4.
���v����_V�C�7Ly�}����U'��M�?2J×j�Ƕ(}���r��Y��L�X
�ߣ���}ꨴ#:+$�Fw�G�;�	�
l��ǯ���
~}3!���l3��HO�D�њGX7��;��յ��� <��#��XY#62�����D_��E�J��k�(�����J��(��f:�z�:�Cn�,;+6z�Q�i�<�.��?��Eo�Y �4ےd"�~�D�o�ŷh�?�lТBX������m�W�:m����z�^�n����d��.�^RYjU,�SXfa4�=�x�í!�Ĉ O�<~r���F��Z�a�B�*��ߜ_�ѿ��-��/�lh�9�.�(+޽�ɔ��}����#m�2R�~"r��m������|a�ຒ]�7=�0Q�C6C�SOy�Az��/x$�·[~	�����,�����]�כ�2K���m(CIS^�+��Sۑ��C���ZP��K�����T�e�!'�ސL�#7X~`w��q��:�X�y�{I�2&M�v&N�˛�,��ʄ���kp�"O^���D�Q�����m�U񼹩o��8���8�_{�T]KrG�T>����4%F�ոϙ�D���U/k|[D�u��(J�*�����:�l�|h���00h~xr��"*M�ʟwqqx��쭍��������E(K�|(j#JER�?z��m��\7T����"�<�a�jm�j�;�S�J5�����y%�^`S1�����������������,7
,~�J���A�>��%�5������c�y&�` ��Z�g�'Ɠh���	�ތ�V���p�`��+`oD�����܃d�}��"����8Z��D��P}{����xB��Q��7�N�g��[ňU޸�3a+`K�`q^.��V�?K��j��{6�U�t����kAJ\@ mZ���/=���1o.�.uA���
������Ba7>��Vmf-)O�+�X��,�����'Hᤚ�b�9[�ȟ?A�2���QfnE�_*�o�q�x)S��F'�cey�ܘ�E�	���ތg8Y�A��Jw((q��<R3=BώE�櫾�>���Ϛ@��%F��w��]�땄QGV��%;--�䥔�G�O4��*UBtp��S�ԧ�Q�g�c���>7ܗb<g��ɍ�����Ƃ���ք�0q!��т��&%���|	�:�q�/�ehXX{���8��$����n���~�\��fթ.j��=�=/$3���-�B��<�lt�'M�����Vf�7�-M_���&���[����;!����u3o���m��_7�
v"�7��aJ�ڡ
�CY�?u���J���x��98z"H_*�HX����Xt���Ta�f����(Xh!}�?����c���O�<��D�z���&rk��j6v�Z�L���;�֫�.O��c��(˧)O�P��Pv-`�j�Q��ݵ�<�e������h>�8���#�,�}ð4|�3Ym��?b�:�gАl�e�Ʀ��R!�Y��J������� S��M��v;;������!2�K6�-��4������/�n[;&�{�' ��VCCc��rQBRq`�����B��!�1�T#��𑜉��U�γ�3��C���k�����g���^���GXc��`�a0��8�:o��ۑ�#f����E������Dl��η���]��u�ip�0��-~9���@��~v�����<�A�'����@]]�E������LZ$�
 �B�|���CC؏�K�d�>lW4��6ţ�KL�-����<"[|��߇�����o�K��PU~���������O.��?�A�v��N6������99r�=���Zux����`���R�q������4��ԏ��gjj��k=t����A2���i�rL��U (/�ġ�8k
����%���Qˈa�����+7���;gg����@�`��5�p�ݙ
�/��+��ԟ�fg�����*�A�q>��/� 3�|��Q4Y��ύ�֨V ����@��S]V�4��
 ����o���ټ��{�O������9DE�te�o#�D���������cc�2��;��}O���������������������/����:����P���q��8�"����K��|,��f���~�'Ic4���#Sԯj9��ߥqo� �\�g��k�F7�7o�(�B� Sr2�cn�ޅ$�g"@M[���������n0��:$""~6��=Z��}��h�����{�	>8JO�]*A xv�(=�p���~hL���#"#?���Z�V�.���ā�ļ�V�7I�{��f��q��(p�/�����0��`�9�����+{��&�Ș܇�-*
!���G�L���ͷ�8�A��^�����f|�R\~�~g�俿P�y(��W��U� ����%뛛�dJxI$�R��g�Y�dX�bZZ�ݑ�������������<=����������EZ�a+}��]�R e����iSԡ�@�Qo 򜳳3��21�f)z���p����$��H"6���!���b��T���|��N����"!]���Mv�M�����AEx���.i��킚ņ탼�fS��3ʷ�LL�e�����O����G�k%��?Wcg��7U���&++�*��mP���%	&�����σ�ͽ�z`Zx:�+X���.<�z��ن�w��2Ʒ
C	����E�^B͚��i*�����Sx�1�s����h��|�Qj�e��)1��H�L��8�"�Y���+{�.��1#�|U�R�Z&��p��n�u�w�j����^6`6Z�1mnӁ���2����H��)@�f@�l��f��'�Jԗ,f���ڤ��냟��P�Έs��7_G����c9��V�Q�K�������J�*�J�$���О�+�G��efF�z��aܥ���$�9��:���U՘�����E��6=n�o+���M��,���+M_1��آ��/�5@y.�۷eh�n!���%s�>�;P+h��ٹj��-��Y�V�=""����2:86/>>>#+K|���?ө]���Z��"6쮝y�^����7�\6OmK��������Z�D��aI-hN�ߎ/������ө�F9P����K�,k��>-y�xP��,/�����G���L�h��hgHZ�7�±�Ӑ}��=5�u?D�G����3�9m-r�=3��C��-ǋ�qT{�W@#��f|�8��� �}�zL��D�:t��a�?��f�cb��������O�Xw�JŞ[pu/[^��=#-FBcҿ��iֳ�p�٦�hT�ت������P�=hoG�V��꧜0�cpHIC�w�� �b�6"��� ��I�L��e��)ڥxe�/��������Z�r1GwHiBr=cf���,�NT�g �����V�~xx8��J]B	["vvv��ё��߿�J@@6�I_G'|k(�N@�����8Ƙ���:��"�w���R܋�Ey�U#�q���Q��B��Q����-�!�`'���M+E�����TR��*�'96�Ʋ��SN��7ym�/�����rW��
�&�r����!-j{qI1!>`��ʡ}=�TT�9�@C�K-�{r�>�I�3�i�a�F���k��;��Wx�_o9�N:J8y�ӌ�rX�7��K���-���Î��^��Fb�������˹r�~u��Bn]H��K��W�+�ӃueY�[���ٔD���0e_�{f93�L�u2I폭O�Xrw �fdP�=�r��%�,�͑��Jn!���TSSÛSטZ�W�$��d��:�ae�2���69K��4�U�f��%����z�#����c%�>�h��f��������z�|����1�e#V�Fݒ���P'���-:��5�ؚ>��d<�^��D��]�gO����,P4��.���*��Cx�eS�,��{�`:{i��r��|��9˖��$gc���@�U߰!�g�����Q���_�+yy�$��j�b!"�:�~4^s�c۪�z��Ք��s8a��k[�+W���[?S+��9����̙l��z^9����� ��{"�]���^�F�x�r����ܻ
&z��͸�P��gñ���W��&o�M�������8W[�B������C����ƻ��D�TT��=<tI#��!R҈4Cw������* (����0� ���C�������Y��p��{�y�����9��q	%��&&���{�t�g,�N�ỰjmF�kL�T����S�5������a	w�Aå�UWW���;����r�_J�!����s���vx�h���1m����7���c_�q�
�͛3��/_�MOGVTl������=��UK���T�d����MХ˩02�.���E`5SqyI\��X����[�G�����z9?�l(�Z;�uL%X�rB���fc�?T��9�<�}���Ltz=gZ�b�����PU�x'�$�����PC��zb�V�)S�"�Fe|6�!~1%L���"+T���I�qis�<����^��Y�S���s���?�!z��l-�5�Y�y��~���<�}	���x�ω�O��=So�T.	-BAA����[K�O.&�XYZ"JJJ�I-,�oa���@dd�sӖ�a�}$\��]3D�8����󍴴�ˍ���ť�ɪs�}�2�m���u�&CFC�ܟ,R �@{��`V����l�M`�m)���������7��߿w�!� CVS���Ѱ��2�L�ǀV�� $ ��w�
U�xB���Q��Q�[���6P;Is�X_�W�]�wg+U��}U+��O	ܜ-:S{Lv_�&�̰�Ӧ;�W&Ɨb�ˆ����k�{LW�U2Z�d�H~�N��l���`��3�bF�J��M�k�ۻ��ł�Ym)Ş7[W��;�uj��l���|���ĝ";���-��0�}����~����iG|�*ˁxr-���x��7�Ar�nyXBB ��H��d8��Z�mk����k
z|Sa�
7�'�����̓���{A-�	�t�=�����{�>�gh3Cșxy��
��n����SOnMALL���J/��U�n��W�B!�o;����C$�n��[fq����Q����r3�֛VؾdW�ן��Ĵ�1u���&�-�uh@D�W�C�}`��QϪ���G�t�g�%Ŀ�f�^����ID�zyx��)�:v"nX�3+nek.��{���zd�h&ɫ]voβ���nY�]�[���L	2�K/��a�����͚� ������@j}/���kѰ�9�`�h�0�����,{��I�]���q��p;_EEExD��R_\^~���9�'L�����eac�fcc#,*�#
ٛ�f8::J�����~�jRK��F���{!+�#L�ä��N��l���<t��l���G�Z44���o��J��Ĵ�U�e�蝿���t��$侧|���^l��疵Rۉ^ߺ��e�Ӑ;��V� ܨ0=� �ո�ױ�U]��gSc��}i9�!3�4*�kdC�~��f���fmF(Ὰ�7=ֵ��$�����>0����Y����;dDJQ�����-dǕb>��ܦ&�Հ���_��`��اOx ��G�5 �l�G;�Bv.8�����S�LA�4�S�Q�KRy�*��cG���og�.�!#ҥ�,��PVn�q<��!�ђ�0�t_�/���k�/Ā}����Xv��Ė�O'�j����:g�!
�����tqA�$�r�D_��533+�Q���F��u!02�6�lJQ�L���N�p����쾋s 1�蕬��'��q>��^Lf���>o��c��&��ݴJ}hx�Lާ�rk�R㦨n ��ԥ��	�p����x9f�稃A�gyݑ���ux��\ݘ6�ϊ�JA���
�z��@���&w��nB9��ʺ�ą��<�����ǹi\*�`x:Y���?��usmw�d	#�_
a����p4|"���G)��v��j�j}�W����\t��z:QM��zFe���X�J4�D�d�=���%�����J}^lo;%fX�Ş�ZD���E�h��YV��H�$�RW�|�V�ud�Sś[��� Ȗ��I�y�á�M���|j{A/�@��W�ߗ �F))�/`���~>J����-�DXZ����je�AƳ��0�.���s��{��]l�����N�13�5:��q�;8����0��%`5 I�B�+�D�o|R
�ʳ�7e¢���g��ߪ���:>9#y��
	)(����fT�_��!�H[��Ӛ/�gQc�C��{�Rj�Fآ���`h]�6���e�
j�ZϧSb%��D�/8%������[�|9���y]DBA(�M�{{h:�zӀf�-�����O5�q����G�C*�l	eee�>�^Eo_�索ۗ���SS���8��h���FFFGs�0���r��)h�jD��$ )��f��}''�D��'�f���@�&!�p��Źx�uu��Ա@���r�-}�o�+Ģ%��Hy�k�����Vx�X#�5�b�O��
�;�׻�U�u�(��6��~`n.s�=���)�A�>6r=�c��VP��H�5����н�{~�E�I�gGlM�B6	�d~�Z��AN������ o�DDG3��Q��]33�Yo<�22(2���%���`�̕�fUSi)������Qy''nM-�ϙ��pq{W�����&_a����`���.->|��)ӥ���<T����n��7���W���4��l��f1���l]�@u���)�Hˑ�g��}_
U�����qU��'��e�ND�Km"I��]�H$�S<��DCE��[�ph\z�i3ܠ�Z��'_��f�=��㩘�c�2*�r��0%U@����/Ǐ��4>��O @O�DRj�D�����.����3��].�������ʰ{_*d��Q�6�O�p;E?:�C�y��!�|�o����ҫ4M����P⠽{���=&�'go
����a�F����'??��xA��������Yyx�a���#���;�uv��Y��Q��<��<�,,h�_9�������W{�љ�ޮl>�3i�{>2҉Yjwf_��Yk0�_X�E�S���F�b7�?���P�֓���š�S�Dl��k�Wu������ާ`��<\��PJ\�9(��L���-�I���l��+w�]4wH��ـ�2���&4��MnB��D���l����;�#	��H�~R�gj/�g�t�};����J~�E��YI�o"۰{;���b�n��1A����/8�������(��|&}���Q<�u��H:�S���s��bX�MM���%�f����vcT�9�J�,,u���
�*0��C�9���s�3�z�h����0tc:�0.������N�?tuj�������M�����c�@��Aޡ��;y�+������L� y;u�W�}��i"�_uo|n���hT>&y˷�?�rk�+èxX�jѠ�6�Y����^��{��ebFH�y���j������nL �~'��V��
*\����X�ݖ|�Cxˢv�/�[��dv!H�PN��QL}p8u
�(��M��P��D<� Ǵ�eF���;V�J��O	8�{��~D^ϣ+Y��z7a�OA6MoUK5u�r�^0&}�k%��} �x[E��JwE�E�K� �����$�<F�\B��O�	d������b���_��(���\B��6�S��=v�O�oju�KE3W+���K:!�����%%'P'1Ȝ���� ��tsg�;�vH�#�'`kף��6J�g0I�xAq<��)��&	<4��i�����~�6m�c2m,����uȕ�\�5�E��I�\Z�\�b�Q�[Q��ҵ����q�=c ڬY;%�K�DT�ʻTmt^���A�7 ��ڶ���}h��g�5�ލGEE[]�]M�jR. ���ġz�z�9���!Iс�GQV�2���qqE�N��%G���c���mk>|�o����̢�Q�z6�^8ly�
��E-��}��?�8���ћ8V��	�-&qV,�Idޤ���G����Ҙ�v-����M��$`��Z�Tk\:z���q����a��HB��'�����U�,�X��j�Uu�ڿ+�3/�lg���2i%�^�e�8�n	��¹�@Q�Z��Iz-}6j�	:*�f.��
��H����r��Un��<=�Xu�S�4h��4���T�K�T�W���K��:4�'�R&��֛9T���#Fp=�Wz+�E��V���@c��[$�O��ԠT�R���=�Z/�Nr�w����9������σ�I�7t+�cp֐�>R4|\�lzKO���C��~�����������-2��������Z���{�.^{<�k�$�~��g�L���{�?3��6I4]�Վ��5�w����?\F�)Р{L]9���P��=ߌ��wl�:y��y^��l�l �y^�X�(���p��z�O�������q1G4*��<J���b��E�W���H�����\+
�5�xNm^(��{�GZ���s��}�n�ڛ��_@Xv�#N����0��ؗE�������VmL�߮E?!��rJ\��D�:MV�SX�2$�ä�����ۙ,�nSǹ�$�sJȑ���ctT���h05���+��p8S~$�"��s�h���L9�v�ˇ�����d2J*
4����$#��C�E�DK1B��J���[�έ">qT|�Zv�����|뿫)��5���d�Tޚ=AG7q~0Q\`_RKu�B'�ԫM�wM=�-�u��/�I����EOV���<�`�gg�*T|Ϫ�������;���F�M
���l���nɮ�P@�H�1,���r�l���p?���Dё&�˝����OVbw[�>��E�Gw)j�aٜ���E9��aU��U��ݠ�Yy��MT���h���{���i-��ir�D���/�]IT�̿�;�+����Ef�����5ݷ�ə�@���_�P5�
���ǿ000�,9�n�v��� E5Wm��p�H)�j���H�k��I�Gg�@��������N$>���$N�H���/A�q��@0z��������	�v@�+-\\��_Mf�y�{N�4�����=���]W���ލ��B�����t>$�� L��S���� R.�Dῧ<8��O��X����ft�Q�����~9�w9�-�=0e��9���P���lu8��y���m��?g�M�% �(��Ti���pt�h��1O��2fEA�<���LB1�c�O�[�F�o��r�HC�z4_���w�e|b"}V"_�h�	�~��	B`WJ楘bN������}������4���Lɻ�ը��i�N?�� Gy��Y�A)\'�����4��D�^X���Ƣ8k!��
9θ{�ʹ'�.w^�����Mk����?��9W�]��8,���?m�<a2Z�4u޺=f������o�)�~ <�����Y�N������:y:�L���;���q�� �u�bc����ȏ����4Ϸ64449�΋�f�9Ӽ/�uo\a�p�T��8���΋��8p��.{���;��V�!4���D�}w�|���p"�ވE��ĭ|�i��e�u �{*2��=��0H����e�j@��S�>s �6'K��F؅6�%�5A>��;�)كL~��:�b}]y�g- nS]�b��j����Pà����2ݥ(����d|v6���n��jX��K�˲���z�$���&Q���Bw�7>�1d����b㽿���������� &��h�r!+q��teP���Z�&�q��t�i�WL,>@w�f]X�O�����c�`(���I'��4�_��1�,���x����-�'x�_����JYO+p;r ���؄.E�Q� ���J�2�F4�f��A;��M;��K���40t���w��Z���?���;.<1+�o�q������Ne;���&�݄���W��k���SAn�I	Ҳpd����*DC6�����+0�઒Ř��&�a�����Y�`q��W@�����`���Ï�|��&���g���T��P'Y��@�=�~*�!C�b�r��^+���"���q��@*�}��e�����^̭�Jd������Ir��n��YN����{g	�����/Ͼ����gk<S6�T�셩�3��J=ǉ�G�iv�n8�Q�@g��Y(?�^XXh��v�X����Ǩ�8��=��Ҳ��y
B�I8jE��ׁS��.���Z�����U���)��e�2���^'K"��p3E�;E@�{�K����`�	5\&�����Yq����L��?h�h+�2���fL`�S��^H�C81Q��w4����x��PBs�cJe�6����`T��a������8�_;��8v��z�@���%�2���w���7Z(`W<@Q�;X��3����"�J }���&���6��7��#��*Pִ]Z���b��>W�k�*���`��;��o�y��b�whŦ��V��S.I٬I�ʓ��� $h����b��R����X<�9-K���4�<�7�����di�9�s0N/�,m0ueDDD��o����a�R�p�"��Ңu!U�Шi�h��� �>NU���^~�C�,*ﳧ����j(L��K��c���~SO�����i $����>�� ߖT��2��@w��<�T����(�� /��i=�VP��ޞ�y�"����Ͽ �&5��0b\T#3qſG��boV��¾xIW�{4�����:V} k��V>�H���w߱�=�i �AWdb�wa�<p��Kz{�Ҵ��t������V	l��!�!����sL%��p[!%0!��$L���W��/j��k�J^�Z���UL2G˱y3tx�z�v~�a�2����E�$��i/�3��#ꙺP�0L��*|hC���URB�/r=���ƀ�-�]X`sj������m�0�@�&y��	��������o�ʯ�e��5�/�H���{қz" �a�� %h� -��:��Cj�ΟgIJ����L�߮�
E��"�\n͖o�n��W"�*łg�cz��9��O�0�ʏ{�:�Ʈ��r��e�@�y��T�%� Mu��:,V4�CVE��_�Q�	W�~���!����E	���O�%R2缢@��*M������B`���[��1<(e�hD�������y����j�}=�yl6���|J<%�- }�TA'fȍ��a!|B�(�+��A7#�^�]�5����ހ�9��K� �v(�kBc[Ի*�_�F��&N�u�����q�w��A/ ?��������2�`i@� ����`^�c������L�O�n�x,��f�V�Bb�	H��?�w��O��#�+�Tp�8%��_U ��`�V�a�B��[�f�D�X���PưD�Ɨ�!�SgF�N��:M���!-�H�%Ox1d+��ׅW�s�=�z���EE��HX�顪���:�޺������k���.��f���G�B�ĩvA�>�o.|o�µ_Qy��dK}�_4��k U_@ОʠR%㵳豣͌
�TPv��|%<mp�w�*�WHGq��Tn��D��j���b��8���ߔ�XA�����X�yږ�kx,h�}n}��dX�ې��f�<��?Ru�};��Aw�[zq�s�䡶d�Y��)�Έj��� �����败+ʀv�N�pAHO�����'�ɚCd�-�V�0����~��?W�8d����Gd������-��Ά�]�]�d��K�b6���x�;��>2��Q����X����di��Ux��zK1F�%"�a�6���!3�";��`��2RH���!yB"��6��2�]j����Zެg{��1j�d�:��J�5	�g��)�Vu����&2�rw[\~�����u����Ah�v�j�z8��G�g{���J�q��	�B�&�����D.Q/��/RV|P�^*��;�^"��	�Y\�j"��]��x��9j�D�c�2F�	�WY��[���k�!Z�5kL�	P�#�<����<�� #���"M�"wAaB�����UVT�b�e9kg�	�E�K�����~O޸4�w2�����#13��+[y� ,&|�.�a���������+��	W�
+*�F���N��(LR�����\������0��,�dGH�\��
!��#Z*W�%o{��u)]V�Y8�b��@	���e��.���a�n�+B+ ������M9Qo�F��&5ayoP�����h�9�F=��%���젧�����Z� J\�+�l��b�w���;��']z/�n`�Si����F�o�;~�P`*0�z��T�F������@ aoߪ��hR��b�����{g�64�A�O9�Q䊞����~z�ݲ��ȃh�a��-u3׉�탛#h`�QF�H�$��V�(�A�I~(�y}e �	��e/������G'�1�i�w$�Aޙ`��M'�phI�|�[:z{%;[l>���|_n�$q�A	(2]f�	�	(�de��.�k���#UK7�*�O�"b��J�JdN�E|�,fog�T9gt�#��QV�0�����J	c�ij�]g����׮��'� �e�H$�R%8X���r����&N(���帐΂x�3/���֞$q��S���� �9�t΅�9��b�e���0�;ի��v�&��CޥO��%��Eϼ�g]n{����G�s�k����U�e_���'b�������́�*���Y٩c`��yI��ߡ �}ˋ�A������u��{�w��QT�:R�P�
#ټ�S�Jm��L�=f������&�H)~�Z����C�̉'e� �	|?��\��H)d_�����"i�i\��?����K}��!��t��;�'��Z�Kt��1BLzq� xl'\X]�T�.0/�B���8=��h��oaZ?&��O��������aL�|���{������jO�+n�Y�j3"����$qO�ջq���a��1)�ƕ ��?�
���s�x�V �{om�ʴ2�u���0ȗ�	���Z�Z��9�&9�j�m%�MAWD_�_�x~��eu ��雹	dWD�����5Ư2��U��A�o� �a�*�Y9�l��堐�e�!o*N#�M2���-k
�����)���A�7�%�`�ƥ0�����O
;l��ЛӁ��+&�����0Y����g\F2uu |w;��o��S~�8�#z�/3:�\nB���h�%5|x|��:����1�ͺ��o��/zr!����6�tZP��o%�]my�xHX�Q1�.��]ڨAD5���[L�_�cYB7����q���"
b��c�9���f���J����f�{����@�&J�!6��	EN�(��"��d3�KU0��0C�O����@u�5�|[+	�m��%?uy��4,d-�����굻�E�I�̀d�]���sv��Cc~'�r��d�;�Se�m�V�2����+�߹릣������(*�s��o�qѢ�f�]��z���O��s��	�/<��
�f7�9��[�:��nT-���;�ǰ'���v]C�?��gV����Q����RO�Ώ�50��B|��$,Α��}H���eu1.�"���FJ���K>3���B�.fr�o�=�*���j��S��	\�G�檳f�[Q����&?�9�o���nv�ߣ�f�\Y��[��w<v3,��ba�:)��90{���H�����"�r�:Dl�1�(4�(:b��������q/aӖ���t�`z��RG�:�]p����4/%�+�U 1� 4�O��0>���H{��M�qs�֬p^���c)VFנ�%#�9�����1�䴧]�v]����L������9ͦ9�������9@�*lo�M�ӄ������Ɗej�`6�O&.�E��3^R�n��0�� u�Ȗ��C��bo���P��m�u��sǧO���K����.m�U>ɋ:�ϼtĩ�k��˯�������Fo��]��P �)�uw"Wp���i�H{�󰕬&�դĶ䳙@JM�vv6�M�8\~8�O�c��\<eX�6��s9�lkKiI�ɾ��Ԏ�y�wJ�^���9�69.���o(f�Z��-O9x�\����]�##���}?=Ɓ���:���L����rfm�x�7` �ʔ����-7|�M*0�{�yR,˔�g��p�-�R̳�=���}^zJE��M=p(XY��(l'��Q�c��F�B�1*���֘��kN;JVU0��Y���kwB�7���-F�3��	z�k�i��U����(��B>�\�Ǉ� b�"o��c�����7��eVd�C��`��p\�9X�ݮ����K�&l1�Y�U'�b;�L���z<�3�t5����iᠢJ� �r�_^"o5��`w���Y��ܬ9t�C���i�����<��aci�����9ϑ�R`<�B��A���wbWco�Mva��wJ>�	]��N�떷#�͚iM�� �$�eZ�*�o���}�W�ۜ~���7Z,<X��Ȕ����`�I���N����$q�B�mbN��ÒI� ���_���5�"1.�gMQب��T%:�֋�Z3,'�UAl���f��|�\b������<5�|�Jw�j/y1����#[bxk�(��=�$� m3��A�D�����Up�3�ݛ���t0�8JeT�^8����GK$;0�s���a�G��,���N�����415"�uM;!(4bR�I2�6_cS�M���f�?�E�^�H����n��y�&I�]g�&'կ@���/h�afD�*rӝ9%k���C�ψN�{��nh�y��ui2��T��s���C*B'�ۙmjy�z�1ǸW�7�-���r��T�z]q��	'y$?�w�}�r�t��x�b����q�}cҔ5C�0>�Y�HjeQ�G�g��&UM�?!z���ԧ܊�`o��޸���l�T��F�Ee8w�={�6n�����&�9�9S'���w)�������&,�{���{��g��C&�(to�Y�:���._��o�,P`�GƂ��N���82�dm����sl���*9:B��|mC���ΒWu�bb�/�K�-,�X���p�ֈ��m��;#pls4Y��k����>��w���ӟ��z�Z<�\7�ĠG���2T��lk�[��/��(O�����PS�yt��B���?���d0�M1�0w���g�4���h��Na��ħH���b�#��R�K��? ɒ����1�މ�0��BP����$.Mܑ�t�%;P ��`ثj�R�b��)�����q<��-�n���^Jv>��<ϒ��ǩ<:�,�N�l�$-�;��y~���vx�!�1��1�q�.ûT���}�O dڊ�QQ�	�8=�{�읇�lwi�kTc2�/��j0��%���ݱ;���bp�h� ��Qx2i�&���1u=��Ty͖FY�"z��/r�{���~�`D�F���I���N�\�A0z_�N1'���p��$AH�>l�c#�7a���4�)�G�{H�拋˱U3�mg/ꃹ�7�]�e<�Q�Y�D�W�#��8����d0L�m/[���V9}�y:<5[����+s��e5�C�}�[��}�_��U�FҢԀP��A<��4)s���������,�`�̫W ���G�	�fqM���%.��0%�\|-r�A�1`1���W�%���I�M��兺Sd-��#z:�%&��c�Gl������>���������#n��K�;�����xg��ɣ��-;��@��ı"v�
���^*���e�����pVT�D�,Y���E����CLa��y�[Ňi�^��G߇���*�-M�V��}o�߲E�K� �!ů�6�_\��-~�拳fq�0�uUK�ԋ�'Ǖ.k�Y�k�p�n�'&x��L���S����*ns�	7%�ؾ��.˂���D]-��%��A7b�u��=Brt�Xn k%Z���zО�ΟF�~�������hg����;�ASc����7���]�#�&ɇ����c��x�BJ�a��׍������'1���,��i��HF���BM�f�3��T�����p^��.�L=T�I0I_�����,��'��B�y��fa��jLh�4ˣӂP� ���N��'�	��[��
cs<��h�%z.kd���sM��a*db�.C|�����(��j>����%�^�,���
���Tt{	V*mkse���<����H�b��Ao�n����뛱f�7�:�u�g)��$��
���
�C<��ꃶ��T*������ �\ ��8��������s�s�����k?]�>u�AWT$ʩE�XJrH�i$�?��,E$,��n÷���ҧ{-*2��l\A�b��#s�^�݇q�e�ɇ�����0~=��b���O#BYُ2�O�䖣@j���	7�/�A4�R@��6�H��|M����6��^�ͪBd��O�z��F>��%��)L[l
Ή�e":L�4�6a������@V���1��c��xj���fRV�4��ߠ�=-�Tk;��>��-pYY"
��[����N4D��It� )s���洒�T�:첍�J��*S�	��}���H.E_N�n���	_N��iɛ�͐�"���,T��w>�i���Ǿ7�rn˖릠��;yp(޵[Wo5~��j�2G�����:/�)��@�+���.��t���I�J4#*+.暇�������Y�w���k��%�J{m�_̎�l�A`���TJD"s�5���w�$�$����������9�u�R� G���P?MSV�2�����@1y^�O�^�m�#%jb��(U�0��Zӽ��@ [�f��'Vd��U�K�b(i�Ҭ�i����e�h���0k�~�;'���O�@��C�]��M*�%�.�&!,��"����Y!�(�����3���T�1�ƞl���T<?�l��v�K&]\�fLK+3��Z>�Eξ�1��bhqK;�%�G�w��K{��r�ʗ�APEg���hC(��B�@�c�*���Q)�`�G'[����q�(0R��MV����XD�Q���|�C��~G�5����Q,#a��å�x�Pd-�6k��!�.��H�]����(%�Ñ���:��v�s����h�x� d95�NM���\!b.�|a��G�uҁ'���%'��U��`�f5Oe�N�}������6ᗓ����k�K��>�����6������� [[!���٢�;�G+_0��&� ���1=z�`�gZ�Vbn�ӕ�Ԡ�o�=sb8[1�/�
�N2�������Ue�q+sB�d���V����u���W�S��}�;cG{#k	`��T<�߆upj�턞�R�#S:P�H�/�?H��n~�[h)ġ��k��4`Wt��{G�q���|�^���稄�5��ѷk�LO�)��"0����.&w�^5!�w�\�	�e͍��T� X1Lr�D�cӈ�Gb_���oߎ��������밋�|C��#�>��;��եE_t�MU�JŲ�%3d�H���Y7��d��%�$_썈�����|����)�bo�h(���;�
������NK���- g�юX�dŶ��Jy��w��f.nn�s��tN}������@�wv����7� �l]��ژ]{:��
uz�\J>�>wa��G���-=_.�)^�opZo�P�#��Sv�F�!�o.0������&f7��@���mą�������k���Κ%� �DeǄQ���S�CX�̢��K�I���O�H��(�ޡ��� %���x����q���|i��	 � ,a:��H�{:������0}yQ�yZ�	�-�]����7V���mF��Yb�?�q:��_��M��:a�-r��M�?���q5�%�'�b��pѹ�
~^nRwwwU�6�z8�m�㱳�Q����y���BK�Y�eD0X�-�6?��u��a�"v!��]�4cز`o�V1�f�����T����&Xv,�
��~�*�.SJ�[V| ������\��>�SX;��kRFq��>�� �K���+Nk`ф��m&�lߗ`�F�X��Q���d�7.�/'�	�L�7��*��q$f�l�>�G�%KI�}kL8�h�y>�|l���~�����py����n{�`M!��5����cj�&{ߑ$z�F���t��ė{�v�n:��C}�[^���}��&+�63Lv� ׄРl�H ���Z"�ۅymԬ��K~��tw�ed&anе�G�;>��ǰ٨I)ŷ�o���/����">-�~_\���J��eYh�5"й<�ԩΥ�
)I�|Ez�қ�X���K>�D�"ʥ���}-�����;��g	Yk�`
��xA1Th�~�W9�r����{{e�&���A��bmYB�# �"����z�@E1�5��ap��r��9k��+�@�P�����IW�N�ث;B~�T&s�i���>nZ�n`�L9}����i|����(Rҭ��A�)�FN"Z�1=?1ZA�q�xF!���K�(��GDEe�#j?���H���5�GCl@(r��Y� �I����r��ݕ����v�ce�"��y�	3�r�ah�Q����R(ؠ ��o�6��&9��w����u蝜fD�|��<7%0Siֹv���6�-��ff��H%zV|_�mt��0[�q���9eBX��h*�h�0�r̘KI��BT�����Xe����{���4�2*|����RyU�/-���.k���`�.#
�-��f�;A���O9��z�5�6�'�!l/��f�^)G�'�F������`��cu'IF��j21�u^[�.��,��	��'�RR|��t�Nu�z�y��`K�%�p�7�'x-+��8���9㍮-�OJIs-P+���wm�h�H���4ǠMq����t���e���J^��5������ud���e��n��/��]�'R�J�DI�E<>XP/(v}t��p�~\�?�o�c�� ߜ�Z�X��)�)ɧ��ӗ��D�c̥X|�jA�o�ܔz�rPHq�ݶ�~-ύ_�/�C��Jt�'9���T1�=[�ѐ�.ū��.b�AdF
�֛�пT%��o���&k��-vi�)vr�-:
�N�s	{ν?�d�>���>5������ {�Ė�_���Y�".����-�s�Ar�XϹ�XmA���Ҹt���)�ж�s^�s5 �|�o(|��k���M{���8�/�&�y]�py�ȥE��$�n����6ی�T$�o����w�%�U�a�L����DO����}��۽��	�1���Q��"�`zލ%���՜ӊ��	��Yܐx��?[�y���mKA߆�dL;�6#��
*�Pn���/s��`�S�m��_M����V��@�,z�V{.����r��u��p!~a�얕��hE��z�)��.���OxG�.g�C�/�b�����F�Q~��ڬD|������i� ���A����!�2j�k�	b�6D��3�7r�֫�j�Ք��R��t.�M&)�4�+����-R�#Ď�a�z��ӻ�{[��P�/�v�[!ç����,m��E������t���"����#��=�`��ۘ��=Q��盳�Bl9�-i	� Yr�%���$��y^f�������q��S��b��dy�	}����5����Gw���j7Q��T�O�.�����p��T�y�Bdc���u�"������̛OdnB�N@���싙
�EH��B��:,u	�`��iVc��ɾ�WϾ�����~ܷ#�7��&�� 6jSa`#�M	�
ˮ���^۾��TQ@:��ě��.�_�J�cN��ޓQ0�H�>����*e��˹m�i륇ia��Ħw��� �FM����H����|��G�)+�r7�>�Ү+�&��T�6���s�4��x��n�ױ�L$^O݌��ux��<����N<P3�����t܈/����� זO���5A(���uzƹU\�Dɚ�X��=�2"��~2}�6TV������[�	�ƌsb�k6W����-�M.(���R�j�wCt9��	J�*.�÷��}O�"�8�K_�ms0&Sr�^�n�@D�����W=h�U(��)�s�Ӈn~2�+Q�� ����}���� �ֽE���K68�T���1�_�����pJ�)���9�D��<~\\�V0��1���&+�w��Z��[���Ǜ͹j+ׁ��1S�?���=��ǽ�og̊�9ԡTU?���-�'���eM��x�F��=�{���sCJ���q �i�}�����Z���li��oY�D���1�a5Ǣg^g\IT}�C�Ջ�H�F������]���,���i����/��s�������k$���1�~pĝ�+ޝZ�^Ŭ�l@QKD�&7�N�x û��o��f{�SS4#���K_�ǳ�5��f��(�x�4�Z�"cm,:����F����"=�����Q����1^��7⧾�����pr����	��
�=�N����˂˸�k��ݱ��� nK�8�~��+�*vX�S�����5���E�*6�H���Қ���煔4*���Z�@\��'��Ƙ�i�����uVYś#:��e�)�&/>j�@䔂"�,UD�.��H]��c|�C-n���%*�tj�U�An��6SKչ����p�q���d\����4���B�u�C*&ߑ`������kv����8�- %*.�n���h�ʰ����S:DA��iiDZ��Z���A�i�s����%��g����u�}ufΙ�����|�~���e�^V�q�����K�gޗ�/KH#ǁU��K̋�%)�T�����zΪp�Sr�f�g+✲NX���;��f��#1���Y�dPBd>��Q�?���Y��Ql�Cu���ޮ$vl�Uj8A.����������h�P.��8����|2'l�{��Ƈ���m��Z�)=�l�$�`�°�q?[�5l��Ҹ�]��EW����j�̺D�̜Z�Eh��~d��&�]t.\���3Q�U��E/������l�|�=¿�����9�ո�Q���uT���t7+ƼW�/Z1�֑krh��??�`�����CYWc���t�g?_����7\���kЇlMf]l�G����9*�\�Рƌ�ǎ��C;R^9>_$���6G˼�=���Q�g���V �E 5�B���:�X�;�21jA}�$�B�J^�T� ~w-� ��%��s#�_?u�;���9NK�j@�(U� �}�4����x�"7�(,�T@ĭ$=��$��t�>nO�C^�m[�����R�SQae�t�dQ0m
|��(%#bh�>0W^��@�suYT(��6�	[3Cj׍Jx\��G��ãڤ�����D��a͝��2u~��vI�<B��6���0Ş�)�g��|�8y&�P��K���C$fΥ�ї��p�4��KC�����Ix ���h�80e���ЎP��z$�q	�%��)'7�������Z�������Ĳ���|� ��_�v�G��FSǿ�����K���%#y�*~�˵q���У���C*�ǂ�L<r�.��8K�c,�+O�gBZ0�O��gr7���9ə�h��I��=m0R�ٱ���v�Q�l
�<�-���U%yyy<HU�]yO�����|6rkE�y%0��L�/b2�E˫C��/^}6�K�2v�͐Wg����w���U��E�ڴ���*�:=(X�ډ�Q,ݐ�}�Y��>�r萦#ra��Tb�d0�d>��#}.�&j�᥀|�MF�,���� _N�CHH�
/fW�c�7	�߼������2�?x���@z��32���ƚӅ~FQ�|�+[1����ݲ�?����O���M}�V��c�e���#WQ��2{S�?
�h⦅ �<("ʷ�*�E#S�,^xXS�tUvc�M�q�|����@H}�����x���L�8��&����G�����IK���6�U�-��џ��u�4��V�����E�a�Z�-5�0��]����\�`{!{!�UC/y�u�����T����Ϥ�0m�>x)X�ԇu�	�b�
 �B�o��6Jx_�r�= ��5��ļ>�����)84�G�xGMr��@�G�Z��E�C�X��ԑ�Ԧ&�E)7kW)�Es��O_N&�ܧ �ՐY��M'W��x��EI+�%C��`D\T�w#|�S���V�l��_�7�%`\��h�h}g�-�DFC���Ʒ!-��D��Sy���ݺ��F��#7�ߩ9�\���AF���� ��h�5u���,m叚0Ym�v"��
'E��.c��[��G_dbF��e��b��9h�i��H�������l��M�gl합���#��}��D��������#h��W���5����+E�T��$��錺�?��֞O.W$��_�KJ2Yx?�դ��R��]��h9���Q�hm�}q��v�U檥����W��7vI�/8;���0�����]7߆S�%G�Ք@�)T�a��h!l�w�J[`�����7��@������W�cۨg���
�hX�|�>ײ��W�!3	�@C/]���PUF_:�KVS�	X١���Ax�R�~��yJ�HA����_�@��i�a�(�.�����<M=bi� �έ���m����@c��������ԡ`ܐ�f?���b����	6'�r'p+��l=�ڴ2Ѫ:����r�E����@�kk�ݺ׍f�'c錒��>�������I��m0�*��d*b� �U���O�=����m|���%��d�����I%n,[V��T��~h�5G>\f,~~[@�t"Ɉ�s��\e�����ᴤh�vUa	�]1& �"x'\S�Y�0�]��o�/�ޛlK�	��	���A�ehy���%�J���E	V�*RnŌ%I2�>%k�@+&�i�͚|���Z��ְ��F6t�G�U
ظ1�;�V���:�cn1�[�qm����f��W��t�,KC."��|�N�,����5����q�Ör��z`�?�ä�Y����[q���o�3��5�NB��9�1�y(�6�-09��8c�S�>����Ĩ��]@�X*��,�Jס.F��S�I�D�Dr�v��:+�}�_�(5\�K+��k���jM���O8�H;'45.�o���Z&��Y�f�F$�R��Op�[�--���$���N��s�<ˬ��1i=pџA��F0���wEG�1�v�{���Z�N����ٸlޱ�A�����(Z�_q�����q����Z�G��]��:t.����r��rׁ�����,���oF���������C~3��,�l��CA�80{�F~�05X|��9�Ϝd�:�Ŏ�5��9��Q����m���u��L9��-�(	wj�}e�-oq�~����H�;ra����?3(�-�ErDz����cs�`޺UU.������ӕ#��5��'�n�+�����μ��뭭>��O���;�[�/�t9Omuڞ��E"3O�^������R[iG��+���_w���?"�����,��Y Y�=��*Q��'�	c/�����0�/��{͟[�r1�Y[��{Lx� �#�� �l	M7��i��nB�w��~���8uM�g������B��8�8�Mm��o`��JU�.�R�d�՜�!3%l�_�|o��p{]��܄\.�4�=�@D-X�p���w��b�ee����""���p�@���(D�����E�]�w#1����fX�fn�*���v��[P���]j�c c���kFI�h��	�)EtKK��u������� �/*�/Ym��el�2/k.���.P'�H'f���*K���	Wŏ?[�������k��vғI��j�7��(��L5HM�,L���ݘ�Y�V�7^c���D4g�t5��>�y�zd���/��&���z��	@���2��A@���-3/zm\��d�@��P���d�>����,A7��"j�I���+E�ח�T���Z�5+'��[�Ț�%M�{���߭p���2~/����3��)"B����r�k[�u��N/or��*���|�ݥ��?d�Z�K�Lg	�8����6�g�g@[��rE��� �#�^�6�@�]��Q��teP��(�T_���r$e'q�č5\5F����N2���)�{釠�&�$�b�.B�E�d�65��;Oȼ��I#H�%r��ڰy�U{��>|co�~^�z��N� ��>}�Y�kQvD�d^� ۿ~�/���~uh?��i������wD�[#�h�ˋMR�糐�`��Q������e�~�,�_*�s�}m���'�$�y���X� �n��KC�z1�R	�_������;� &al�dvRb�5���A���c���
dd#FA�A0�+����/�T(OӠ?���X	���Ҁ%o��Y6�eV�����5�]���]��tl�X�:.������[pM*H���Ӎ�����N�tk��6���rp�̿�T.���6�x���9���k6{u7��ǡ*|i#Kr�G��Aæ��K=��yynl���h6*��#�p�VrT�Z�Ɉ*��`n��０԰�ɤ���Y01b�aY!�b-�c�����B���2V9"C�m�y��,�MP��˓ǌ�}壻��i��<}Y~i�9j�+޾`^T�g��g����EW���
�`|����P�p(���D���툭�Υ�Ug9��f�{D����㥺�w��v���xn�_y�N�$(\.RFNO���d@����t�}����Ȓe��ۮ�a���W�oPPЫ�/z�~�5H��X�"�UE�fC��  J~<#��UP5�q����y�Z��D�yF0s�����"(�c��$Z�(�8|{����:����� ��u��#�	�Zc@�J�v���7�8b���GzxE�N5�j�q�GD��;"@U�����W������oe���w�y�`J@0ȋ�� ���8Kz�\F�kR�.E6^��Ś��6f|�nc�e�ۛ����y�5@D���LÇaDa��ƍ�A�Gl﷤���U���N�_���rV?���r���@����F~Ɣ�e�K��"��ƞ��sO,*��J�Аhb����#�i��f$����rW�0����E����N
(�-֯���\[py�R����3R`_���6�xxˣ�њ���/���WN$gf��X�� C�t����_�z���qu�ݪӼ�c���P����R9�w�o7Jf��$�$����8e���u,�b
V�|� %��8E�'�AZ_8+�*��v�*o��ϒf�]�QA�T'K�P��w����JO��*��<dw �z*#������Π� ���KvUL��v��p�V�j6���D*��3�����w�m������=F�s$��ʱ�-pu�@ٛcMm���]�����trJ
��sWlN/vx�u��)f�3�r[�{W�N,׾f�v�"7�i6�j�{A��F?_�1\�ש=�w"n!otFg����p���Í��_�$�A<��ԅ�.�' �\��,']T�+#Uѻ5ɢ0�b:�� �����o�GŅ�T��v��u� �.��z���>j����Sd�՚:�e�v�WAś����NI#?<�?7���M�wH��j�cn���İZ5`�����aۂ��PO}Z�4T�a���6�I�w���^�NC�m�Pi���4S���i3�85:v��>v#;�s��^I|�2��Wg��H���/�������<T��,\᜻�q��\�M R���S�-t�L�g.I\Uy绱���w)ZL�v>B����D$q����ZĮ����90gԼfTq��k��������)y���B��@��xL��w�F��� 8	#.������$k#&����k��lP3�)�ڈ\�d<�����0��F�s6�����d���vʖZ�*1�ݷƏC���a�:|*muyO�L�zO}!����莂��(�=�g��i�����Yy?~�i�4s����$a��$������f�^%����r�m�A�u�zP�A�v�hm51��}=�MM�u�C�v���_)D}��v�B�rߩp;�RM��;.S�:��w����Y�+�Z�̺��[�w�F��Y�)`�h��`�P$��9�ܸDѼ9�K˼+*����XZhĪ���[Ggq�l��4�]���'7sT�]�ѿ  �8 ��@���=h%��RLxL�˸��K���贕�wL���`}�:=���'Q���a�����5��>c�.�z�8�!bd7���K��RRf�w�!>�$��R�眬�9"����Y7�IY�����[�mo�R�q�O���qZ�6�1md/�L@���SW��H��La��M.��Ჴa�vݻ̈́'�E@���&?��;q�T�&L�kp�B���:�5�x�|���ٌ<#˛>�����ٙ.S����[�!B��~1%O �����v$0g~�|O��5���$�!�xi�+S*cEY=��H�V���v3d���;��t�-c��$}����7ֻ=җ�a�p��p'��it)��8����{�)EE���/��63Xz>�]�h�4~����69.��G�ά �+���j�q ���Tr�*�\��&}GZ9N"��g6󔱣٭c����n�]?ρ�+G`���Z��K�ƭ?�Z�m�T4]L)Է6�ye���*[1/�_n�Dqox�.J:�[��h���D��%)
PQT��:���44���0���{��$���J1��%ѥ�T�S�L/�V����� �NY�Kv�s����:�W��{6P�W>�����dB�k�j6A^ճd"8g�C�t�h���J%�:��qMEc�c.u�%��r�2Vw��m��n�bAمX�:��g9'�r ��O�d���=(�\���y4�/�K�ꌌ�n�\W��A�Qe�v�G�����+@������l^�ww/���1�T�3�{L�d�Aʧ���$��l�-�Wc��T�/-�9�W�{�7P^B�Qv�>����zo��h\����{���`}�(���}=\���n��� \ɿ�Wd����*HW�w�y+�K�V���]�G��t��������������v�䫁�e}`�(�#�՛qa|�o-%�"���i@�D�o�ѿ�g￙K���&��MF�����4V �ti&�ٽ�J�m���V�!�~7B�$H�^��9���}#�L�A���`ձ�t���#�дf�����E�s� k�|`�m�!�Ljz�T���d�Lb���P~�;}�s)�g�o�kj������L���W�����ё�zňF�.�_���a���IR�����B}�Fy�0p�-� �5	@�A�]���
�^����M�D��(L��A��O/ā�#D����k%�ˢ= 4;�������n�(�.Z����Y�[�)�M�˺Rs�E>gK���j,�):Ϡ�ʕ�F�X|ҷtv&��>ֽ��x�h%���S��׏����܋=$g���=�����n��%��~�%�h�=	��r�sX�|p�<(Zsu�0��!^-����h��OZU؂�Y��6K���~�7~�s"=�o3�e#�FJ[c�^2�8�1�n�X� "T�L�%��8-t"���k<�������x�M�N���G����rV�űa��h��hg޲�/���\H�v��/�1�u���e��P�c��0��⻣aagO�ׂ���^�O#���Ay�y����;J��s��/��&� #J��(m��MJ~"����dUm*�@mha��-U������1�a�rz�L��I5!@�r �y�ɉ\a��l��n#�:|zߵ�"B�"*��U=�{����K��a��Fu~�2�Tml�j�~Q��Я��v����_U��Oۆ)`t��Xpf�U<����*G����1�$��Ln�v�5nTE�G���� �>(��.�	-8���h�1m��y䊖����Kt���=.��&���.+�z�Cd�Т��p$�>����V��x� �-��<U�|��/@�n�,�ݖ�W��o���/=g�%���hy�󶳧�"Mp�ꍇф]��!��^�梹N6
�|����M��5�o�ni1��=�g�mbPZvvTFiV����WO t�f��$�l9�I�XY��7���ޠ��5�lK?�˫ّ���~�9��V�����}.�(�ש���&ד��l�Stn�V0P`PG:P�����>�V틽�ۣ�����}1���6d��T��:�?�V�:����^�����r-�%\LT��J`�:��v_U��D��\�=�����.S�\V�#�\Z�<f�f�1����ԩ$�y������ �z@Z�NU�{Z@~'�?���tY��;�-ʏ������4Q���y}�IX���Wۆ�&����U��*��^�r��fV�����"�Opkw�BU��vo�\f���w�͵�����ޞ?Z�(�{p�ae;6��N�� B����97��S�_<��1��V��� ��C���×Bmu�822S����w�<��$g�T���g��*�9��>���mK1AZ����(�ޡ��_��[g��(�5� o�@������$ҡ6�A�ψQ*I&+�0r���Q�Яl�}q�}n#�Z=�e�Nq4����,��@�x�a��]�&+�]���h��u��^�v�z�P��o���H��{!w��P�q�I�rs�<���>��� �@�y�g��4Vt���zC�Fq3����Q��l݆̍�0y?�ډ��Qs��f+�ᔳ�tH�}��T���P��K�'�;�ks�{�#~�e�;�gT�p�WVW<E�Eg
)S��^�P�/�'b'v��o�G�;���+�"ك�B)&8����r~ӿ݂���6�!�Lc�?�%�4���B0��đ���	)G��lܚ�n��R��ͳa?]��ܫ\gjp��
�:�@��S�����v0�Q'�o��sȟs�uo�Ћ�G�@T�^�b��*���D
P���}�S�7q�}� �#_Q�>C.�c,]�}~ɷd�.x�* ��q � �o�qcNm����7?�gǦ�Kce�D���{�4�\�F��&;F���_��~_�Q�.���r&�	d��8q
�D���:���>����bB�N?��P�!��� t�?��W�q��*J����Sĳ9���Mb����d���j�[�ɱ��˱��pKg[��c�
g�!�Ѷ߀�B�@� e�Zu�Y���2&܅4l���t��9��M�l��2/ NU�w*��bD�NC�#�4��a�/�����"@(Ա_�5�c���2�����N悖�3���B�9��-՗]�4�P��\���R��{�S�<Mw �ت��H-��e��+cɬ�1M:��|��������=�6�Yp��}mrr4q�����E=L�Yr�L!h
U,�0"�"�%��5=��T��y�
���`����Vi�?@<���ϸ�Ρ ݹ��_\_W�ŭpp �4z��qc�$�V��{�/��zZ�9�F��C�g)r��^r&'|l���&�fg;��T����]�GJJZ|�)~)u �!|��p����H!�i*f���6v�uI�����GH^]z.��o����wMP�l�nq\}Y'�d�v��\�I�4���t�k�7L��Q�%��NޓtЯ�V���TO���#��P�a0�u�3XC�?�1�z�P�q&ZZq�� ���o�571|A��Pq|JM+��7|_CG�d%��ZW:��.��ȡ�\yu=0���7u�!OGx���פ�+�w�F�i����CB�z�8�ٱU"�k���a~A��Ўxa-��s�j�(��%hTu����v����H��X%��G~L9����U�*/��+����>�$�r7��b��"@�#�����	�L���k�7����,�A4xT���"H$K�<���r�y� k���r�1B��h�H����/R-R��[éݱgL�BtH��:|�+�fNG�嗾"܃AY�CĲ᫸HX@c�f�6,�"#�i2��ɂ���NF)|'t�^M�.ُ�,����B���4Э)ӎ��g�o�>@[�'y{-�K�!���:*�EgԷ�(g:��X/�>l����{A �8^R���bԗQK�1��^^��N&⽝_���\�\@�1˖,v�$�S5#\���R���0�}�<��\�TJ�����o���"�HkԞ����0rb���\Å�a7��2c���悔2������Fp%��Ϗ��1c3>/6,,��A҈�￷�"�F.t�P38N:h��`��ॿ��;����rTπ��=}Z;�h��p�q�v{}�r�{2��p�ҜU��w������, /�xqD��@a,�֓�w@��-0�<w��h�;��BК��Q<)q>EU9�r��%�E�;�pa�����>jo�Ǒ�ڣU6�FJ���V����'��8g�#�J���|�c�k'�]Dl�|=�7���3:�!QfU��#���^O��f,˩��A>���MI�b�v��ڑ���jxz|~��q��6`�G�˚=~㭙�����~��Kg;�&��.�{A��\��7*��n_;�	�Ϋ��Gwm��鯘���X��y�wa��P����.v��6�D��aX�QK��Ƹ��n2�j��`s2C�ޓ��O���e�*�ngֶ/�]�-�;��ot �h� �R*�c������*Ⳓ,�GV��=�¶0l3ih��dWG�Ð��V���y��#tV�Um\��	�Uh�0�3��?�jgFx��0h��J�$s����P6V�pkM^_� �a^a����P�CS�Y�q� x��~Z�$��4e@&�j���F5�2�����Z����U�'@	��� f(a#9 W�)�Dh���<'4��B�Z�b����CK��k-�O�pg�۞� &c6ȭ�Z���=u���)���s��O�~�=����?���['d��,�y�Z�t�:抣i'n�t�e���.� 9�uS�%�>-��Ce'y̮��8��B�A<���t;N��D�bL�4�����
��0��KU�w����[Y�W���A`��w�"�����T��_�+�\uX�8G��T�J$���b�~U�@yNc�%������Md���.��;�>�>�s�������w����,݊��[�0����2�d������չC�V�AM��������,O�Å���Me�^�>���*	*��-+iG�e��} S�(�]kh`0�����%@B�Z��]63����Qp`��
�a#=�)�*{צF��t�7/�Ѳ_�����b�I}mA+�{�h_�CɩP���m�:�YG�w������ŵV"�1��zA��a~��U�)��ߢ2��H��H�]��LV������0�V�����f�us�!���j���:�@^��,df��k0r�?���� ��p��r#[8�/m�s�X�VD�p�$	+���ԹY�?�c�&R����2m�o���Ƈ8�\o�ޗ��L�Җ��=t8�p��O�99D��k�	���o�^ӏ�t�>��e�����}�䦫R�}�?���_h �0C�~g��s�j3��`'�N�-�GD�g��V�a)�dj� ����0ᰴ!�#8a�������g�� ���H�\\�Pn���X�"�+ a�j��`uyuu��i����{-�d�)w�h�_=�+����5iK�y�"����ܑ��#�x��pr��W(��2�	T�Fx�:zf(6���V��ܫ�Ta(�G<Y�&�l�kc
�ѝ����y��D�n�����h#�t��Chճ���q���u������%�i'�	@5��!5�ڹT+g�+yⱟ���U���ӷP�7Uڒ|�MR����Wp��S\#TFIn퇿^�:�q�w�F���\��h���<��6�I�d0���;¦?�Хx��y�s��Ua���ay2<����%a_V%�tF7|Ә���t���(@�Y~2�8��%]���A\;��
�����/_��|�� X�D[-$A22�D�J��U��]�����"f��}S��(��6�$CSa<�d5gZG��_}fe�8�3��v�X/�
K�U��'Z�@(@{
�����_հ�	���<������ԭ�� �c�Qn�������|�ư`.���[���4���B�&������`���|"��oa1��$|�=�<��ִ��+�]ʥS#���YDP�bcC�܆�ˏ�� �l�BӶאF'�g#7F�[�+z��hJM��Xx��Wv����%��9X2|ٕhKp���+Q�q�e�xT�{��̡X���A���}y�M�UY�
���UMp�":Zuw��,z(٥���p��17��#�(�,�-����03,&���xx��
�����<�l��ё�3�{ٟJ����hd���ʯ�{d-xU}�ћm	�c{n��K��m��q���
�f�]�n� J�W_�P
��n�$����<L�ͱ�	�u�Hz^u;�C���	�/b����:�sCy�'��?h�'�Fy�� ����sQ��k)�qs�?�_?8}Op�Qt���I1Z�;HNIy�j �VO���94q��s��|5Sa�Ȍx�Ɔ��Q�>�q���Q��N(����������.z]h3d�R|����"铳%p����G�����8���0xG�����#ȃ�S��}y{ ��.؁?�M\�UƎ��!����a\�VA`�>4
��Ȇ+Y&��;�K��p��^��&�ggx��\e?�c�{H*�ۮ�أ:ۈʧ��1W��a{ۜ���:{h�/V'�� �:���:�x�$�ȟ��X΢�~3�T\��}�xϜ�`!w�����u$�+山����?i���Ok�q!c�����E�஡'����=��=t@�O�b���&%Y4Z-j�F>�E��ac##@�7l��2p*����T�CE����W/-bq��d����פq����V���&]|���/�@eL��E���n�J��2���#]U�hE`қ�ͷ�ē�N�"JF��<���P���(��$tkf�rf]�>B�3ag��t����4@��qxk�@�:*
ܼGx�צ&�$�"�S��ֵ��2]��9!�����A�`���[�pa�H�:/��<�$*&�6���y0_k��
�=3�u�w�f���i_[���Hw���:F"���|��3�C�c�X��pg�ecA���+��0�D�`х����X���O��rR�)*�<�|��S�5�P�ְĜ�v��ʕ�GJ��ltΙ�,H��UFO��(��tǬ�5<����++��H�C�T"srh���m9�w�� 5�;��Ї��h�k���#�Sx �FE�ҭ퓾���z�u�WD$�����e���%,88 x�>�~����	�V�!L~�����n7��-��I���zX�M3Z����r�������ut��5������s�j����#a�B�?Ĺ�m�6�QF?%���h�⚠]�W�������u��0>���iz?.Uᗉ���.�+�wJ(�@�}�����u�2�h��6�	�k����p6ʹ^��J���.kon��qk~`�>�G�A
��ƽ�ko�iw�nw��8��]y|	W�p3��ڝd``�^��L[��;��@��&N�/C_el��te���7�|H��ż�=q�14��Fy�{�Ju�����2�5[�W�9Y�}��&��E����L2w�m@�-��RM5A�._�PSR�<LB����(��I�.�8�$���h�U�d%� ����6Y����P���Q��J�;:�:�W�DF�%33~2!e����xSh����M�%�B���5���x��"^�O�+g5_B�M�S1%���9�d�Vv~�/b��C,����ET�b��� �`�9,7�L�\$"�2WʡNZ���I�ᡅ���T��GE�R;�t����a���T�f�H%����#�`s�Y���1|n`j�L:[��vx�7��ad��V�$�r?��mǙw�^���:���	DЁ"Lr�M9��l>r�uO�(U���cv&�c}?C���+&YP�(�ѵC�e�HbH�����J��M��l,|S�&�,M��v�o1�?;���0�{cMU�����@υĒ=0:f2뺗bV�?��������ku��Y�������߸�ʢ����9�6����t̸*��a:�<E���dg����`�IhCk�	ӊ���`��-R&�p&<S���'�S4�ɍ������F8��M��!{FO)2��n�wq�.W�;U���qUI�i�_��3E��Y*o�����h��j5�N'�;�5��4 �:9rB<���,^4,�}hI")-�*Yrj����1p��,���B��b�K�@�g}��.a^R��^��F5%��d���dk-W���B6 �NH��Z��I�,Y�i3�f�Z�u���ߟ�;�K�q}j��$�Y�]�7�]��nN�Ex2RP���Y����	\��[D�9��L��f!^��aY�������K{�ԥ���}����x�{�d�Mt�(�v�@��e#l&<GKDewv�.����60��%��,�F歺�t�'.�}�Ig*�-ג��&�A�w��櫓7���#��]9���'���r.o�5r�}W��z`� Oa��|3	H�6&v�5�ᴼ.(��»᥃��b�����7�@����vPQ��C\ȏ�`�����J�BL�ƺ�p��[
��M���|�Q�òz,m��i�%���v�P�����F���M�H��E5�C��nS���E�W�?�[Մ���{=�n���Zބf[�Z�1б1�"f|��������V</Go[:�^eS��]���*�l�4��&���k
Q˧&R�81B��NX?Y�r�Ϋ��V�F��Oϴ�IB�+{���͜aq�������X-�|�Yf��FR5�|�{�	��O���i#��g��;eB<sV�**G6�/6�
�pf�3��{�
w�·��o�"�Q;���v;�XӂS�x�S���W>��pn'%�@�"���+�n?�����eo�: ;�� ��Hi�~]0'|�`���B���h����@[z{��9��'�k3�֛#�td�&��&?~a;��]�\�zpE:0
��CP�y�fɂU�6A�o�?�7�7+&޷N�*�وƦʝ�i~�l�,��P&k�t�K��D٭�����z !��8�Bʉ�HQ����F�������e���U�3.�G����y��ˬ��Q~)���Z��?*oؚ�z��|�09�{w�T���������U=�Z�����	���	@@���ú��F=�(�I�W��1" ���X�0Q�Q9��i�0����;�RD�����?N�I'���z0a�Kk�0� �OD�~���Ta�M�1O�!��cd&F,��P������#���5���~���qk�����Vg<���<���0�h�e��ӗ���zo����F�Jc���N��W��74��c�Sg���R2��Z�j?ػ��p���9z�6}�ҥDb�]�u,�2x��Yf�+�z�m3��D�2>q�!���wV�Z�X���:m�,�"��P����й��͗PF�K���Է"%�Y.�
�6�P�B�����@|�xM�J��'���0"�VWs=��?���,w���2(*+ϵ���֓۶�I�d�1ҭ����׭�p�\zz����+���9���Ֆ�O�!m�h�G9�p�5P�xT����`$��o2�\�MJrR|u�H2��o����C>'��]�΍K5�\-�̠[�<��0�Y<�Δ����
ysd���ji�!���4��rҕ��K�,/���U�g�	?�L�҅�x�}%Q0�y��\�B!! �`D�6���M����wTN]DxM����n����}�"`�`2�v������X*SGǏS�ܙ��HL�#�a=T�z�#������I&u�����]����ޘ�
�?�����ի��bS6�#ӗ���)vAc�vߦ;N�Υk�.�_���h�U[苭y�h�]�Xq�렟����C���&,�۟�os=� �� ( �{�}�9��Y��� MZ�
o��Ԧ�j��ed��2S\�"f
�(4� �ܰ( �ӻO� ƕh�c<��*~�+��}�/RB�	#������n���{!m!tKxv'u����6��������;�]�u ��#X붼[u@}�_�⩁�:.��?�9Ŗϗ���;�~��pzl�[�u���!i�D�T���=K;mg�X��x-)��`<�څ�x�1�Q�	�1�{&u�H�����7G�9qy <``���\χ]4y�3z*�RG�c�J�XXp1ғ��!�ݲu4�M �?�/�qF߁�ˁ���?�ы&1܃�$1��@� �!���5�n��+}Z��v_$ 0~i�-b��θ�3��gV��~�������-�S�+z�	X4��CR�/8Qb��K�K�xUNإ���=�� PU�Yz�D���� �a�3����ǔ* �4��@���"�7Xd�Q�(�K�R���W����G�O�q� �aY�s�/��^D��t ���{ �����W
D8*������p�k#wwA��cb�6I�tx�`S���8m#���5PD��K	�g�DJ$go�z��+9�{"�BÄ���0��;�,>ļ����[?��� j.�� ���	ڋ.PW�`bĨ-�x4��j:�؇�4�Of��W"�b������Y�������D ���/r���g�G�>ɿ倿��qo����������!wח��O����t�������'��x|H�=;p�{k��v�HeI�{$;�o��`X�|m<���ߥ��l�<u?�t�^4��=�~3\¬u:�����W�Ҥ�޿3�p�j�>�u�oϿ�Jh�f�ʒ|�,N�ܿ���/TK��������-�)��>TK��f�#ѕI�X�KK2>�21ʝ�e(z�E�Ow�RZ*� qeb�X�� ۊ(����.��b���St���"�h{~,���^��/��]�Z}𶀑VZX^B���B]ő�v�o�j���~�����v@V�_�%H϶���n���|l����fC�}R��Y�a;�ϔx�Y� ���h��?�6,���[h�`��V
#�2�㔵y����~;IX�]�22\h��$FpD���xz˰6��k8���݊�;)
(�]��B�J��w�"��C�Bp��%��>߿�G�s��^k�^{�Ӫz�|L)�u<v�*f��wg��$��d?u�B�d�іٗ��C/prr�X2!/CR)q�i�����Nf3�偲��&�9Շr�4̜�h0w�kc��p�����4�9L�y��D�1RD}'��]�;?�.*�{Q�q$�����[p��ѿg��=��s�lנ##���n��;�;R%����[���~�F�M�����%ݷ0e6^��y�8O-1/r��Jܧ�(��O;p���B"�
��٫�.�y���L���� ����e|��7C�필ӈ����9>��W�3�� ��FhV!�&�f.
�ƕ��W�s�	]0x \�å�Sa��b�e��inS��-�Y��$�Q�)�(UMVl��j�o+���TGן+Ƙ����3�8I���m�w�-9�K�{�S��ŗ��N���I޼�C�u�{
:���{:>G9C��o�q�2C������r����Ҍ��W��3 �w��-Ї��i���t�"��X��ķ�'E3$�Ȍ~Sx
;���8���`ec�q�Pkn�d�����񊥪D�i�] �9����!8��5�I��͞�]��wc$TT�\�2����D'5�b$�ߪ`6�`s��"�J��8���-pI�o�J�H�ߏ"���������+1��)Kq��m�Jl�f�L�:��1���5)qZy�Ej�G�6{!���ơ�xs|��s���M�gg��ͩ��X�C�����N�������nuEt��i��J��9��F�Б�>t�_�Vc��RK��U�����o����SP�W):~t'��-ϗk{������.}���M	��a�oR��$xdC# ��n"�&�|L��8�@���Us*��ñ��#�g�=`�x�"��{��]�t�Fm,}�U@��>G��P�rꄴ�$�l*j�8�g��
Sj��%?��獁�Hy/7۾�[�ô��,�U޹ś_��<���p!}pz:��o�4m�����u������M|�T���D��m�����'_iP���(�B%��`'�d���[2�f)be�Y@�ef���D@�Qw7x8�i������O��`S���"������9����:	��$zS��p��=B� �.�,+*��7  �ܮ��>�c�*&(�*F��4�"ΌMwvo}ixkn����T}C��
�F`�5hk�p{ ��0�����: �@ʗS[X��uG���[����h��;;�}�6+�����3s��<�|�,�/��t��bu�����"������I!���T�Z�������xo�)��~�9U�.�ke��_�f��t)��'���'��3ة��߆Y_Ts2K�#��C��k���C�-{q�������"��L��{z����+߶E^�P�<IS��;A��A���{�����������K���P5�6yDڵ�S&�PF�q�_+`6Z�O���W�������tG��<�03/\̰:���Z"d_�M�?s>c�m�]���dx��o�5L�]I�sQ|	��,_|:AC͕������6H��Y�*�5��?�V��h+a�4�V�'n�}��֔�M���u৷A'e_ot7�kN�����me2);5�X�i�3,m&Ry�9�qE�kG��. Di+�-A�m��=Q&�5�a9E��.8�'�Y� �k�だ���0[h��>�n� H}��=��0�8i����?��ǌ�d����"9%��ز2vɳDwW��㩗�)��/3-�uhp��ϷTw�q2�y�H�V�i�����u�����_#���o�&/O�+����W�ؖ6#��n
 W��>	<��)(''QZ*P̐M��KH���K�|��$�A�-*�"�\Pxd�'�����h���7�T����_Q9�ߡ���,o�V Z�r�w|aNw.��b��d�߂<G{lG�{Zqy�2X�껶r�8s YXY�ż�j��7��ǽ��D��/���e�Xۇ�� W�6>��/��a��.��a�B�*E0�v1�H�3Q�x�R�0�'iʥ�dr�S9�	ǧ�}�/kp����ꣀҢ}�h�O}��h���5O����m�ď|���ُ�+���e���9xY�k�#��#�'����nS���N^��L�����)eY�Y7MYmq.̷Ll���{Q0kױ��(�T�*��5  �e��̕�I��1�v�jzuO-��G�<��	�:�u�S�;T�ЮZ�'#�� �R� �6���5X"3'4�3�� 8+r����+ǓT�8��sL�~����6ߟ�%���}9���|G,������?�D�͢;���S���bM��C�i;E5�|���`Jج6+�%:5��o�z�V{f
Ǝ��_�)*J4>��q��3�ʻR�I#} 	뷨�3,B�(��_��Ti��p��|���W�eD�߁���\���Z�O��H�T�*o��?o�<o{/�D��ru{˘1>�|�~�՞ 7�ϼzx��Rҷ���8���F�I�:�O�oe�Rh'n|r8��.�F�H��7�h�?S�����y�
��T,�P뻑lp;]JW�;D�5�U���KFzkL�n�����U���#J�*��V.�O�2�x��-l�������j�o�P�����2��;%@��Ija���o��?0"�ҏ���lCO_����g��_�1�>虝گ�I~�����Dl<���bD�ia.�O�ˏTRk(�OODb��S�,��@�`�Vi�#����kJK��I�DօD���Yt@�l/����� Q�Ճ2O$����
�c��ST;�G��J��?/ 2�̡ǝ*p�̮m1�����c�处�:O��Sq���7$��E���HD����v��Gܼo��"��r�f,�jqu.����}�ؖB��U��+w���g��ᩮ����� rҚe�0� V
��#���e�W3lҩ�4D}���$.ˡB� L��K�8�_�*�?��Z�@� s�WFt#ƌ&R"L��MQ���lݾ��O�M�H�|�]���w� :��]����p�۰ge�u��~=�Ԅ��&�@E�_���������VO����ʬ7(���wpw�����a����'�ܻ�Û�Oo-^N`d��QH�$b&�����Qd�]���K���i�?��}�x�r�'b$���	�Nb!w�W�#��>a�+�����t64:�o�
@O��y�\�s7�}ɖ����:�g���9���:����x����6��g����uSi7��[�~V�'�����l��MhSsN�����+t�H�H�reL�ز�iF�$��e� ܱH�̱�u�%��F�"9�I�E�g�~��8!����� X��7�!zBָA��u�b{:Y��^�qrJ��e����� ���%��.����N���[��'�÷ZS-���7��"�M�����v_�㓑,�[%�7/{$��w�(r'�*V'�y��_���Ƿ����{�Q��K-���\�/5|�K�!���Oy���9>0���hp����v��E	���9ү�i�g�8�e,��&�&��i>q5��$��\0��腙=m������zQw�j��"1�IR�vGY���>�}B"��b���?�"=zM��Ӓ��r�3.�ȴ��<[���B�8]-��*1�ZY=G��+пF����&a���R�f�����o�*���aB�/d��F1���j�z峌�twgtS�^�<P�݆������l|^o8O�G�]d��p7��d@,��	�Ɐ�����F�ʾҹQ#A��KW��հP.��R��򷍌4�MYz�y��TA'2�l0=�-.�/0�K�h������[n���o�-��IA����[�ǖ�c�-�~�� ��x��)�J]���8�R�J�"��hv��0�ۊ4h�b��}�O���0����3>�K�O0��1|��;�Yb���il�F��������C|P��{��,"t�*r�&��"�y��8_����[O�B�d�~��4�m]�>�����<8&|��%����F���L�@6x|�
N��Ic<����UV{�hE�D F��S����G:G���X����aiA�	8#�6M�]�����Ab}�p$���l(���dNl��I����8��;D�<�&��"�g�a�L���%f��|�m�1��hlHQ^�q|��
w[��%���x+yŲn 8�.l{�pyz~���k����[L=��7v�mga^���~����cYo��T��.��?(��M:�K6=8���e���@Ba����m�y�����@6M�����]ch�e��7�鵹�(�nG��G�vs7��_F�n�C��|�:#��D��N�S�Hy�/��n=6��ϰQ,;e��6�Y�w�`QP#ޘ�`�i���Z���/,%�_���HlCi�>�?0�&4>����ƈ��%`��Y��t^i2_�6q{���������k=F���K�����q�y:HMf'�%n�"��
��!�U@ ��s�g�ǲwbC~"E�����O�O<��B(2��"�)��:k �fB:ju�;���-J[{���=&f���D �I��yEҴ�r�~��o�俰�M	 LI?:�8V��LI^b���  �9�(�g�r����MuU���u�/�l<�cb�k�~v6����*�2Q*�mСνg�����w������Ԗ���^�I����bL����i�bΊx���۱�v=��r��~����f;��s�0U8���V4�c��u�9  ��7L��
<O�=���8��?����+� R>V_���`m?۶�jG��6lq���+j9,��0��7�[;�&|+������C��F[�#�<	�.�hA���Td�#����b��l7{��d�.!�I����n�&���	:<YC�y�K�f��ԗ�4�R��G��p�c�g^?m\e��4�$w�SWՖOM�&�<R�k�o�f��i�/�HLR �p�|U$�꿷b7�@j�`�Bqf��A�j����}�7t/5�7�xu�h'��n����<��5�D�N\z��.�{��Q�aS���Ӿ�O8�~�
����'H�9��/`���u�+2�꟎"Z��*L��3��Ol�_�8�"9p񦋳���'"��N �!-j �r1N5QQڅ5��=�N>���ӌ�Gk�J ��
y��#�G�\ ���{�A�k�;>y�Y�?=Z}��>����<\Y���V�O�u�5�r��KF��5�W�T�O���3J�[%2����h��gY��z�;>z���W��&�D�j��yO�H�Ey�XL%�=�i|�����]|�3F�w�z�Tr�z�1��ۧV��d:�N�E�Iǽ��-n$��K�P4�� ��;rziL�U�J�}&�@�+�a�q�Sѿh��=�&�
�ox̍�%PbfM�2�7����As��L�v6(	3� �1�2�)�<( Z��J.�|/�U�ҏw���;�;�t*���~j�G���g�n���LQQ4�}!!�c�t"+�a	��X.z>%�����gu�3���Ԙ��}�oP&*lV��X�s��K����	���A&,i��j�o9Bd���4=������:ZE8�4� {�z���Y�����'����ܯ���L>Ԓ�W���S��k��s����D���l	��ݧ���ICvC�����S�3:WGX`��f��K(�+h�L��=O�*�֮�t����e2�alFi�p���Ȉiu��x��N�?>b
G<�3��oz	xm|��5R`\PXb�D�A�;��D���+�[{�޾?_��n'�͎��!6�_�f7�{�/;(;v��S���q���d�U��(d0e���M/W(���/�I��9�/
7`��o���Ԕz�����R#	Q����7I�����+��G��u�ko�ਹ�S.�x�t�7R7B�s�{�d�R��㾔߾T��c:��;�?��L2չ�
=8���m:�]X���nr��{'�˜ZdT�܈.s׋�!8p	�}�+�.�-����5�k�l�u�yxX�N�����zs"ٱ�9�xGݸ0�tb�U�b�5`Ob�IG QV�J�2{'73#�O������	&5�	���õ���?/�>�3�U�Zl��""���H�aܚ/ �`^Mo��|�TT�e��J��є`C����������!�[�
��;'&���<}�Z�}I�?r���MSF��Q7لw��"PLap�.I�K
3�&Ǽ�]WrjS�B�̎�Gƈ��5{ү�����W��8t�Ө���E��W5��qmq�^�2��@�~�_�CQ;N�N�:�wU�oJ�5���
�g{�NaV?�di��o�x����-a`���!L����� 'úO��Z|��4�i*����Q�f��������ͯ�����3h!Y!�n�価�`�T��G:r8)3P��77�T[0hM-�~��!�� G<��&�4��t�9ݧ.��7��딚܆��0>��wXdP�!k'��ֻ���
Y�]/���Z�,�p�Fk`��JF!�x�",��[cz�V	��0�Pv�ߪX��<��?Y��-�|��FH�}ʅ
0w"� f�P�w�w�=aȘg�\�	�}��`J����ׯ4!&������&w����_�`$������:��4G�}�W�5�'�~`�� �l� $�����4�}���,�h�e�������-�/E��N&BO��)�d�j1��G��ڵ1p�K>�BQ��C��I����F�^3�Q����ڄ �lU�F��X�Y�� ��I�~Z�� `n�z���ӄ���PZ�\�
��z7_�u=L���ӬU���#���i�A�"����c�q ���K����G+���Ujv���	i�������j���.o �M���#�����[��ۏ�G�P��OV�GJ�B��l@�����&g>oNy�I�*�	�N�u&��ud����Y#�jTQ��D��y�>(�X��0oG!����H�>[�� PW]�o�n���Z�
۸zܑ��}���'��J���v��\�$�/ZD�����j�X�ґ��8�m��/RQ�GȲI��V9�l���`ؠB�0][5/edtoX����2����s���	o'���l{������oyl���F�R�N'}�-뵮;���8�'�õ�Ȓ������}�0F���ֽ8r���o_��3^>3g��zl�Y��)��k�Ax˝Տ���ь-�K�(�B�lVv"O�a_}�3�w��v���;�ЈW����������+[�wI�l��6�������l^�.8���'����&!~��n�+�<9��X�+���ߑӀ�n��w��9& nQ���OU[Mě��5@V]y,�p5�k�<�_�Fd�|�o���>�	�1�����������0�}[/Z$�c�'�܀��c �R�Q|FV��ŧ�"y\��P����x�	��FT#��o�R����5GފfǪ�>cGo��6��I�����kBُS02y|ԏ##�d��\c9�zk4�)6�|�f'g{����Uy���ѿ������k�u\6��h}�K+�'5����ny�d��+�j�UIA2������=>� έ������D�V>a���}#�dR��2?�I���j�К|�$�xn���޽!s��C�r5xl���|���1-u�4i"�B��������Pm�n��^����\��/F.@ ><)�	�,���rQ�+�38!5t�p?�Oz�t�b L� >�~���~,^��T��X9����ى�8H�]�*�$�y���A%pѮ����+�OOr�j
��Ta"�&S@IF�/!��j8�4��T���QvCqC��O  (M,f2�g!�,����)֮
��.�Q	��׬���B�	��6n�.i��87"�ɼ�{��;�'��I�3����a���c�V\Ɋ
���Wx4h�n:%+�2O�A�0�!7��Kl�步����Ĵ�+;��xs�!S̖hhie'Q|5�!����b��M#�l)�6c5�]�'|IV�B�h�} �7_*����/o�25̌���E�W�Y��s�GX�� ��<#щ���xy�m�g�]Q%f !��ޤ����Nj��u��H0[�1]�/_�f���6��]��|������!�E���*�*��B�A�@���Q9d�3�t-	���jdHJ��A��zQ&L#7]�{o�@o�%e�Ҷ�~L������SC��vEl�LQx$q�N��zo���7�;n2�GP�����~�z�U�z�}��0-�1Υڂ(�I��Z1�Rd�f��5��(k^|I^0��� n�)O�N�oS�&��4!Ҝ���Iu0��[�o�1O�#
h|���.���:�x��l	�L+ѝ`��d�����*H(~1! F��|G3%ǒ(�\�1t�m~D���A���GJ~Ye�J���D�U�C���أ�n�)^���e��M�o�Hq��{ ���$����'X&-;�(+��E=A�ڀs��S�ll[�*���x$�Z_��k:���WQ�-(����#z�1X�DRk.!|�������\g��@���f��$~��W�k�dte�-i��!��L�����!(�6�j&���MO��P�~L��kdG���NdRcp�zF�^!_�#ᷠm�7�2��ѫT��=��$��앦Fm)�7�%Q��}���w^��Mׯ�V�7p�*�0���Z�u��(��+y׿���yS��#�Ʒ��ᅢXs�0 �m��ih�/`N��eƉ9 |�$�[� �I�dô;�q�2�Z�|�`�]C�tB2�%��&/rPD�4�Y3�K`.�Z:�8vK�`��6[�"�1�#j�o(�N�,��&���s!��� ��d:�nIz��y+W�,��FN5V�Mh���s�����bm�������2�i~����_-����_>���w�䉱jM�:�m�K8�%!���WsIZh�h��ps�Z| ������n��L��?�v��L�ľ�"�$���]Mޘt�2�R��I�%�g����Z���b�������g��A�F/5�Z�Ga�{��
�B��jL��x�ㆍ�=��	����,��q-�)��}�&�7�&d�D[�3�>Bb3�D��%�x�{5}]%�Q�O:��?}�$[���vl�X��7�1��Շ�D��)^)T�㾯4� ���S�Z�=�{���X�x�3����5c���C�4�H=��s�Q��sa�X�9�,L!
PBE\�d4U'����s����Y�p�5Q�� /��>����כvXp�Ł+cD6�;w�zjמ��Ͽ������w(}��۳z�c���c�p-��r����Y��<NL�K����X�N�=y�W�������"��~���0�*���m����ێmy�>����S$l7���oE�~�	:v�0�{y���3���� \��oj���Ѵ����V��}����տ�!�yY��	OJ;o@�ٝ�t�P���o�&oYݸ��o�*=���c,L4q���Qz�1��	Q��jZ�'LkOV��@:6�?l�6�F9��5�
�����b<��v�gԙ�F�6'@����Q���ljM�����?����L�)���N�5�z��n$֐tˤ�!F���mE���2�Rs�vS?�"?L�R����7_f{�DDR�|l$$��pl²�]ICK�m�$���tZ� ?�xt{y�E<+�|�[���,�qy���z������~K��J��4ZE��~�&�xcT��.���#^^Wv`D�QTQ) ��K'H֏����9�2�ϙ0�=���p����dR�\���G&���^JD�7@F ����Ǟ.`%R�����ށ����TN�>�n����{P��͌c	�>�E�m9�15����jz���Е��Vy]z�y$��aw���t�~� ��c߂��M������U�9͟5F��x=k&�4~�3kWpL��Ol���\/����gg�;�g�-{���1��7�?p�A���#���qU1
ݧ]�X�����G>��&����Z���='��C��J�%�rc����B|&x#�����v��xR#|!�25�ֶ\��f��ψ�~I�5�ѡ��`J���s��S@�D1��M��9�݆�2
�Ʉ��G]����Z��Z�:�7J�"W��-X��ʼ4�Ub�{�M���w����׼��#='�J�n>9�/4��1�$�x�6[��C�	{�C�k`4�s�#�J>�'u�}Ts�<=F��;h��i�&�s4���{WSo|�(�Y�[��B*�-��֏5��#��	��l����r��F!���+���F��+ }"��m6���Ó�c�(���R����<K�fv^��h6��J�����clb�"Fu�&�*����(�?�?�w�/�K�On�o�D��,mV'`K��9�2�À���԰=��RĤx9�34��'����K����|��ھ��.��Ľ��W�q�:e����	����Ό�$]�A��]@at?a(��̧gYρp�_�����إ(�X����#����)��� 1���-/�"x���gdc�����U����_�o��Bss�M|N;o��f�ݮE���pA�"�{�x̟�f?]g%K�M�{�N@�D���fq��r����F�#?�
\b{�P\����^ �y�Q��n����.�S���׫ժJ��K�ϰ(�JRX�nOV��p��w�D�^�Ej��Ƣ\�HS�G�'WN|�d�I�z`S4��{ �}�߬l9�+�g��ג& y$S��ˌ������g������C//�������9�j��l�.r���Wb�^����(��aEM��W�)�/Ϣc�Α�iGw�Vi;V�:A�H������D3�n�9/���VsE����˚0m���M����+T���d.3��=���WqN��Ȣ���-��~ �9�Rm ��g;���΁�R��6�Z{�%z��l���अĦ#��Q�֡T��0�+��ðQ+�ڴ�3���5gꩴ�΃p����q\��7\DYi_s��D%��4Hi7b~X��CL���P���_L����i�y��&�U7,s��X=�1d9�,����B��~'��߯�y=Or����gǬ�/j3A�NfZ����t�M�X�G�G ^�פ~Є�Md-�v*$���w6`�/����Ǩ�M���{M�3R(��n'�����u�����̩�z��D�n�	��Ď\]���΄CN8`���,��ǽ�f>M�.Y[�V~5���=ʉ�r��E�-����1>F�2�n脲8���p^��I��wo	�PvI)����Z��4��'\f���R�*��J8�1�k�K�uޣʠ�̩=��mZ6��T�\=���#9��NBbg{����G��D��}�%3>�ˑ�'����]�ꑿXo�v�H�p/�Y�_®4�h�+FSt��_�2�؁��6����*|6���`	�yk�㜪�v|5���T��6H��"|�P�5��{+�D��ѴC�[.���ǹ�U��i�3"T��Л�@�}����e��4
��4�A&K��	�S1\�g�d�@S�$�?�Z$|�	�"%x:��D�t��=8Hj����e?[�[�yu5���@k�Ņ%i� �,�wʏ�ӛ��B0|^r���+��3CKρ�NE;��z�������������P&���/��$A*a�������e�G�eP���
��O6��Q��]gӋ]�����1B ��`[E�&)m�Bj��B1�6Y� _[�R�%`�R���ڏ+�A��҄N �%���WX/u�U�O|�>�D��W��P���t�V%mn�T��=i�3�nJ�+4Ŵg�2;R�?oN��=�"I-�nzÐ1k��aa����?%�]���'61?��ѳ��א��.�^f�x7����L�z�ю�f!�����%��b6��x!�����S����w�����M"�B��ִ�K�ΰ���6B�5�M���.���5D��"ݸ/����Q�V�_a�,��$)�K�Gd6~�2�kRd��Џ�K��Z4�\ئ%����[=���J��ٗ�x(�`K,�}c��3����++����?�|QX�W '�w;�/1���%o��>���w0g��}&٥��a���;�M��ռ���c��I�ڼ7���_*\�p�U�A1�X�X�͟�����y�E�!ͥ��}���1��{�cF;*��<����ʨn��[4G���s�U�{��9��n�<�����abvϼ��}��ɳ�����?NOd>�.Ҙȵ���R�M�]g'�+��q9��r��[� ���|8���݆6jU�<L��C�O0_��H�V=�?�?K�4kF�m�5�F��'���&'��iBY���o�3�;;�u�Z�ژf����;�͒1�f�������;��R�Z�Y��}� ����Ͳ#�A-���嗌r�:���rVT�J�Mb�Tg'o��;e��,��=��W��X�����ǟ�oL0�ʼ.-]��گA�G4���������D	��J !�:j$KV&���p<:��8��{�JVAb������yN�I�AW��.]�z���`����ꣿ��<��x��؁�J��0�|���_�SG�g�C6x}}M�I��i�3�ϱ����әK�a�χ�|�ه��	�/� ���Gf�W�{�sx�糊�r|��\�ڀ��'s�F����"x�z���y���y�����4�O�3
mf�;?�������ۧz�-�]�_�#Q�n~�ں�����Tzޱ���BN�ͩ�S��?g|w��[}}�Si�R���,��7a�BA��n#ɶ02���_�S�35ܠ�򚟏�G��M%��1�NX
�U�`�!��SC ��\Tx#1�]:� L�	���'�tO|�����V������l���!@���M��S[=�TR������A����"�`M����O����\L2��h�P�.3��n�zw2]�����3O��;GZ�ІS�Ǣw�7�CT���P���}[��ֿۗ��#�6d�ĭc���
0�r/�������;��ZK��OaQ&\�;B�֪��ټڍ�G��?e�"�3�g\��IN�<'z߲���m�<�xM�ץE�/�j2GLt+��^%|wd���2h��^4G�9�B�����ɥ*��9��ۭ�˷�BQ�!�2�F]��?�O}#�A�֎�%o���≦�C#d��q"`��+���^t����f��YLX �����'�<O������;������_5�!vy� ��#ոG����V��� JߑqD�݊���^R��	.�����4R��V^���y!������;w�*���z�&?�s dY��,��n�*��o�W�O1�����E[�`����j��6�&ƫ��C�nY)!V��zDV��u	���.��9���-sV��(��?Ƥ3,�o� `�x2�P�Ki<`����E�]��-�\
�Qk���&��s�/F���&$�M��'���w��eV!@�l��b(�2O�.]�6p9��dc�W����u��9�
=ū�it��8ĝ�!3]�ب�̹R:.�������V+t��-+]���E���ʪ��N��{PV���@�^�%\�m0w^sn�$V�N�|I�7J�s��´|o���Â����^�>��f��-���3�7���%�.}FϿr2g^����bz�2��� ��6��DDoW=��s��c����������Y#��
�G�3@/Ϸ�O���+?M�e֩6,�!�0�S��G"������T��+���[I/Bc_�ne��#3�����Q3&�f�H�dk|��F4�އ_�,YN�w%���V-3�;�B�W��R5�eECjw�&¤���N}z�mGJfT����̿�(ޙ:ı[�
' x^8���H22"%����ˁ����wy�75�F+#����BY���3+3.*Yt$EYB�1����v�+�W���I�6J�9E/�p�!�'a\����a��A/n��u	������q�/1�ӄB���[�,R����8�~T�$�=�!O;�
�\��-�M+LK��I�����g}�[��R3h����x���j�$#dIͽ�-Bų\�g����n����'x�=udX>�f�3��:J�����[�uc������c�p��⓹�#���[9&3�W�<���&R�5t��̬��t���
���徚��:}��A����@�C�;U�2�Ђ��0����L*0Fϯ��Aq�T�y�td� �,�eQ#���[|(��L�d+I�[���
܆��ITd͋��D�Gĸ͋�����gZ���M����8������/��f��n�����v�[��v�w�|����
:�(���YymO�D�#�ܦs0�����~�s8O���u�~e�q�1����Ru����*~�Z
��[����4��bc����<f頙�P�Ȑ�C����,�``�(G*5���>�[j`� ���O�ái�=!3�e�%�Ж�:O6��-�3��!��g�����Gi狏�09�¶���~_N
9�\-��9��A ��1��{1P����	iM7�<1U3 ���KB���[�.8��4n%x�_]yT��'�i���7^u�ҿ��!�4`�U�K�38!�W7/�䷪Ӟ��]���V�p���K[=ـo�S�x�{7�[��	^C�{���:����gE�P�g��!��{�У����:����U� �������'`�<~�{�9��E�P��0�~+RX���ʣ���[�AxQL�����8f�ɷ�mؐ��j�4��
�eٴ�l�qW�5 �Ʈ��t��L*L����u�%C��Rm���Ҿ8���������U&�\NU�B�D��L��P}�4L�i7r���S�R��MJ�]s���q��z���}-�|���	�������p2_ռ�A�[]EdQa�l$�mngKu�]ns�w["���~Q�=�-���0|�|���Q��L��H�M~|�jH�谍W�(5�M���U(�X�ƐA���U��0�-���r��ve��Ւ�aMo���u�U07����Y��P��~9�ߍ� �>�`t;A��&� ����β���O@8�b�H�l��b�F~��J��~��ō�������Q&釙D��k�ӗT����s8~�UDT�`Te�&Q�.�ܼH��-}��z���kp3�����0.:��9�2sA�O]�}T�y�H:�� 眄I�v|c��H�tլg�#D�TM��u�j%�o�[�6��	��Ž=1;M�!˸+��"y��F��-j��*�#k��dK&[��%��$L\��5�"Ԙx,��H�ԋ�:'?8�v�'�
�3�7yNI5�=�y\�RcYIu�y�����+t_�;�pF�y��р�c��$NZ�^��`�j� ���������S�ݙ�o��ܸ����ά,�e�tt�l�����v��:�$y䲏�\�]� {����$-U��#���K���]�	��*�`�4��̘�ALS�'\��*�gӵH=�¸ �R��T.i�Ky�o���U�gE����[�����bEoD���fM�^�:���zķ��X��i^��_'�??s$-A}��UbA5��sZ�	n���M��8�?ڿ�	���)�����伢�<�4�~�?%n�m�A�Ռ���mIp"{��?_iX��
�9�T�WP?��l�՟6��,��"�B�X�$2ޚ)�rX��K��
9b�8�4*��7�ޯ��aYݠl0'/���Z�&;��Q�q84��ؠFԡ�2��%�7c���PZ�LQ<o�r�?� K�� �|0U�������lu^U(e?x�ժJ�A#Jd��>�<I<A������I_����1�M��N�HiU%�$@9#�T��o��.`S��NN�f����,;��tM��>�s��u�ͺ'��I+q��Z;Uï�K���G37=��e�m��AAK��U�[ך�r�����~fw[�e5Ӏ���}Zjվ��&�r�{>S䀭��n�Xg�'R�����^�N%�dԞ��F5H�_4 �q��d�ܒh�8�O�+"
�F(\�;�I�ˉ�ooo�jXt��t{�W�/0	�߲�y$��~����M��)Aj�59 ?j���z~��T
E:��]KtF~W�cR�[& �F����M�9?��K¿$�,j��.3����5�QI4	��ZWݥ�b�$[.aP�pv�J;�D܅�����8At�*����Tޝ��sG������X������9�IB�	����R4F/Lr;��������C�"���ʳ��3<a�r;MG���v#q*pO@K�|�/�+N>>��:nc��y���a__��<I��A�ʆIp�S<�V��Q�7��\	݋<� �^qd.]���x�2/��I��౞���ިq���� �5>z�X���y֍�O���Н�������	�|���n�]����N�@�����www��.��f�{�[�,`8�twU�]��Jf1�����jB�]Ȃ�1���d^m���R9����h�:l����zd�#$��Ɲ"O�/��	�Ï�g���$�۔]˃B�Z,�K�\�ޛ��z=�~�����-����y�G���r�#�᳽f�������V�wI/7c��YQ�rr#�ۯ���s�S��%��~��j�2BK�������*�_���w�w�63���F8f��V��t��8�����P�;���$�R���>@�E�H)M���|���q�v�v@���[����c�G����s/4��-�,1U�����$/X42r>��M�����)�<�����h8_}]��4n	?�&:@'J~�Э�;�eç3;=*�H�wM�]	�tѻ�sB}ͨKK�U|���vh"��2x>^���"^��j�q�c�դU?wӘɎ"O�]��-�Q��=�����ѡ�R=��~��1��ܼV�������:�K��\�%�z+
"����n�:UI˼g�\`n��LTO�Ŭ��e �<�5/YYT�u18���UF\d�>�=�����9g���x���۷�xR�D ��o��n+@,��05B9�U���<\<��gB���o�}�A�b����ݼ֣�No
(�Ե��޼�qM'��镹�>��]�s�TY\�O	&0X��|;�`>!����+z�߼TWɂ���W�Wӱ"j)SE��0o�Ku�!���B}ܧ;!��a�5*��xێ�>"�;�<aO?��v؜��K�[GR�ЛM\C�+O�v�0��b׹B�a�`�4��,ܹ�	��Ҙ�Q�*�;�(�z����(����F�����C.YN-��z�dy8���Ll"��6]վ�d��7�~R����z�:~-��z�ID����c��_�Sy�����S(<~��
 �(��}M�V�K���-���{;A�T�N���f�xGP�k����J�����ͼ�����J��;yR��,�B�;~j�0km4�l����JG���	�y�Ds���k�?�
7�H�u�TI�Г��j��b����(���LQ^��+�F2\9O��l�1S_�c���툎"R��,�����2A�}xv����䝻�O���¨�^dI�4�����|5�F0���U��]d��:����	����0h�=h��eY�_�q_��̄���L��ĺ��	���!�q�ʓ�V����+a�űx�_�)��)�
d��QLN�"YDt��,E�֧�be[���~������3���-Q��/ߊo��D�'$�)f����	t�^�z{}O���wT�=7i�K�>∕��5�b��49�F'�pr�a$J��oEp�Z;u��h?3�kH0��Z X9�G'����)I�8�,��<��]����r��������B����6)��A��G涧�9� '�y(�/i^�S�A��G��u� m,Иm��=�g����a��K�h>g&���8<c�4�,��3�^�CN*)�n)1�3��ټ�� �Э}l���4�[�9v��ֈ�1���=H`,)&��\8��q��|7v�g�{�JK��K����V�4���@�%�g�5C�	~�i1�j��4�.�ok�b��9�0����0��4�#P$?j�9��pF<��l�!���חu���j�z�߷)C[a�d!�1����}3�l��O���r&�<+�c�����d$	��my	0 	z�[昬okk;8?�����r��P�������ء�u���z�3��<vi8�n���H�o?�Q
��>zbG=�L�q<_�v��&q�q��!����9�V<����v�1ת�{}�ԏ;d#�'��3�4�@�6w*d�a�agK���R-�텢����d��g"������O�÷i��Q����
h��^b_<'l�;}W��3��Ry���3:Oc��и�%ڜ���5��HS���n���ۗ�q�S(����k}=���M	�[����sE�F�[#��~�QlD�1��C���Y���[%�o�RĂ�4�Y��+]���=Q���:�:Yh�?��e��[N��(�'5��(��G*V�s,�l���j� ���*.����:�=�j/�>���o��{��:���?�g�3����m��|Bf*TG�Ԥp��}��8F��Q�w�	E���$�d��yP�S�Z�
������_�o��W���k��C��qT��?- **j Y(4+`�Z�D۹��}eJ��9��9k���A�f]O����TQ�勾v��G����B%���g՟Dni�#�d��BX�Km\�3�s����lo�T���v����3����6V4���m~Q%��-.�'���~Y��]�֛�l�Ӓ�S7�xZ���,��d�w!��U[w�����@���->��<���RRs�V&p���zȜ����u�4[>���9*O���R\��(m���ڈ�(j��~�9�ܙ9qy�B���?���9�����U�f.@�a٨���m+�2AAAw��Hk��������*��o+�d���v���ϝ��L��_չ���B�5���z����9xB���xpԷ���LoK��'(鮴NG˰EĻ_2HD�8q1[�"��H��5�\l��@��7I
܋ۍu�{�g��6�ǟ/�顿4:��D#Ժ�x7�&�(WKF��Ğ儞��Z�뼸�����K�#�Tm4�����staT� ryr���Լ"v���9���Q
Ţx���G����-������.<�w!�=��@*zT���k�iE�.����?���������-��@.�Ջ�����t�nP���r;���}�yjm�����z>r@�����_tn[C��O)K��g��6����d*0�V577;,Ynn�c��Z�`�!P�_]�plC[���@N�Sa:�q�)�r��ssy��_���c0�	���|��bx4�02��r�2T�nS���>o��h�_�6����s���ϛ��!�E�t4)��&�G������2��#�Ay�qi�=�����8�JF�n����ֶe�|F�4�"X���	f��n�!�0��_X��
�ڟ��Jʛ��\�g���}���=J+�*���@:�s%̍����Yq�Qi|��A/`Z�8f�N[�<�7���Z��é'yCpp�r��P�dm��'�7ukyB��l���N^���gn��Y4K;!
�Y���rqsA΍<-vW"�'''�����`����dM�ű���ӛmW����K�� ס�� ��EA���˹ž��C�����lhB��~y*���r���zSx���tؔ�v��}� �{{�hw��[怰XV�Jʋ�b�w����?x2�-Yu�!���{I|��~�?
{#�zb ��4{������l9kFYn��h��[DjX��ac[����a�6K���h3^�O2����烠�ȋ]!C����Sd�b�9 ;>������eZ[�3.�w6�\����p?�����^�q�C�������j q�?l�A�u�3������J�ݞġ��Ђz�'����r��5���{�*���U����$T��� !�;Ef'�m.� *0�N��+g,E�S����;6����R,du����to�A��0��w�\��\\��t�[���6ś`rӎ+�U~"�~h
����)�}�->��
pޅ��љ��E���!���n+�Į���<�����m=��q'�$����R�ö%��3�C�i�$����}�p�2�s�O�zy��"s��� N��Ӕd���g �}&�L/����*��"!*����?����p�F9&ggM�W�r.m�re�NjX�fff����; Z�Wx��\p���(/T�H�E~��z��]$���p�n�^?j�
�~��������c�v�;�Y���+tf��kq��}H�!�h��(�H�4��\�����%ǯ�����='����P���o��j �!l�?�tːʹ���	`��vl6���T�������A
��oX9��a&hEma��)L���0M�#wY����C�i�i�e'���ƽ����!W���h�6�E�S8;W���QS?;�n�:��jD-y��/r�76e\��4^^q�(o�R�N���S9%[��vl}<*q��պL[F�y1����@���*����7��oB�:]�G��) ����3�x1 ���Q�znz0�Ie�^%���J�(�ງ&�M���ْ;q�^K�w�ζ�+V˃N�a�-Q��w�2b���N	��L�d!��ąnɉ�hҡ���bd.�e���ƥ](�~�n�E���H�fiV-��tT�u��ψ"C/1�齊�]����,8T�۞#�ፎ���=����r���(>�B�{4���ͩ;Ù>ِ)�)x�!�P�B;<x�=����^�A��BT������àm@*0ğ/b'":����Z��g���Й�Q��hr�P_�E���y�B�N"8�:�%r_W����|܆���Ї�!W��BF��.�����Q��Of���|h&w�m5C��p&w�_�p���#�2~���:��O`�Ԍ���r���K�Ha�ז�N W��4b�d��-����b)o�E"sV[0<��'gz�8[i�_2ljU���C7t��~��|���i�/��a���p5������Fi�� nj59ԠE��#?c��J#�6N�6�Rƒ�'s�o��X01��t\H`d���"�ٿ��Uf�kl�!BX�����ܿ�S��UA�V���^�MWW�9P�%���B˵`�_n���tO�Ӷ��:�_����|�j�01����#s9�6~oo�2>c:I`�o� �ɄH�|61
��߅	��4�y�����\�C������-��k���ٶ�L���}��6[�M�z&Z/_���%t�2P�LP��b�/k�b�9�Ţ�^��F���i�v�0�XC�~f.]���m�Rh�$��8���uϘ�z8T>�k}ﻄ#Q��$�w�4�TF��ǌԽmy�v�R� ���\�:�acccm����0L������鸑zd��۶Q�fG ��4�"�i���{�@�n_LlJ8�2R�&CS��"u��Ö��t�X+��
��� 
Z�����,��v��r���NJM����1��&�0X�n"pђ�����|��*�+f����_&�m�L-�?�e�}Myq:-���-Ow��}ኵ�Q���IkSG[8�`���Q�i���F2��l�8Up����r[�(��Q�Ǒ�w��v+��iI��B�o8��0�?�� ������I)��[�V���d�abSp��
T�I�}Ӄ�F0�c*%c����Ҹ�˅��;	/3I ��=�D7\�A��?'�/��mK����me���&e"�7ʉ��h� e��r2��v^�$�0'Gf�2 p�6�,��ez�P���1I
��i�1g��:kA�<K |�W� �F�D�6�J�@����9�����=�N���������z&h�Y�����Q�����n�[8�~96�~Z�`$@�qy����>��h�ݪ4���
�Z�{2��W�!Ui��|xl%~JY�g��}4$�~h�M�s�%��@��L�*A8���8�^φ�d��
�����J�����
M�$�$ ���YR|���N{G��`��-Q���`Z��o��kSO�EN���z��`错�%����RH3
�����H'�2�L\���TSC<��'!�/�QĠHקa�oEd?�>=y�����佝��2�J�`3�bS�T:rTDh��	Q0���i���<ĩeտ��a��;%!B�!A�WYL���?��e�8���}���P���Gdѳ�m������4��{����E�����U�~BP�f�5G��用L��G�3������u�SY���Ͷ��˹u���$�v��6�Q�`i�0���]�U���2�hr5(�b�"Z�^��]H
qI�\V�����ûu����J$
�������H��ƞ�x@ҕ��/N
�a0gu�RӼ��7�20ۥ�j��O�v�U#Q���ۇM��u��̴�5�5t̝b��𘜙�|�>æMt&y�Bh�;�x*�r���D�Uh�YEM^�i
r��\�]\T�V��S(�şt���<�T��8�IU�,V���@1.�{q�7n�[����(`�އjq_ �^U�J(�h+�wu��ۏ���7��J�F�.�%��VZ�EMS\�Jd3���W��7����9YI�'I3��"I�,�C�$��z"�&��SsB�nߣx��IW�K5�M�GT�nmʯ҉��Ө%�C�9����,)l��!3�:�՜*X��?�U3��À�qIJ;n�?\�Ux�I�|cm���ϛ<
6�,2a���G���������a��h鋡������Y��G�`O��.��@�}��x�|���$Y�GlniAI% �s�/hH�R�#�j�sȴE����!��tLF^���IU���.���={h����+���%��Ă�HX���7P��-�YRkB�f"���w�c�¢�\�V��
F ��BIw��d @Fi̥��6�;=�Q���ɏ̒C[� $N��YK~�h���vbp�k�����ץg��2�V��a��U��&���U�k��+��v��Pv�l(����S�P����<��Ce��6���z���"W��͋�}#�B�ъ��a�+����F�Y,�Tt�ܩ�yr��
��W7 �m�gM+�}Lx�0�H
x�<���+���y&�gz~�2��Տ��C@	��O�����C������K')E;<���M���_vZ��MxU��S��u�p_U�n����M�M��2l,��9c�P��j3�|�":W��(z�;!���,s
��ٺ�:�M�]�,��32Xϗ�⭟XNd���Vx�i�e�[�8{�*���;4+�]�ŕ]������4#3P*���t�{�zs�q��Cnw�$f6����}���W������\�r���GS%�ixEqȢX��Ey��,����!Ry� �`�#%J�����cŢ/�J8�����9e���F"��G�谘z���Fc� r�����x����
�s����gXj\ઉ��r���>1���ܩ���S�@��E�ف��o�~����f�d D)��l�5+��۾ �ߦ:���nnn62�ֺ��/��񢀉��-���|�.���`�㹲�f�c�㲆ow'��gna>�׀���0
{�An5iW�����Y�ɏ'�:{pb�����������N�{�n8��#j���2�&��-9�0MLJ%��I~`��:W��(�/ ��e�TUgKu�-`Ђ��@��V���1k�k]Ɂ6�.\��Q��DC>@p��߿�節��tnu���Ȓ~-Iֻ2�G��u���g&u���RV���C�ͥgLi��h�F[�:� �%�ʪ���2��'��eaF�l��~]�����ϯ�b�nn��(��n�	�'<Y���P3�H&�0�!a�,�zҎ����!��_�wϢ���o�9hH)+&ѥ�
"0���OA��^�?!�w���F�5��|�͑jo��DT��q8��p;5�����M!�r �I|���z�� l֜"�������.[6����~��sop���С�~:�=��	𐖖J5��顈��	�D�wL�Kkiiu�8����>4?���l�!���-��s2�"
��ݩP9�/�!nA�j��a����ڔ���ͯ�#,�!�0�Bg���8�����aS��\ %�~NY����CJϋI|(�B���׍�Q~t1X�M�-��p��5�֯1Ɲ�z�͞�&�����RXd��:�A�Y�-B��̺ף�nޟ������ED����G�u~�(ذ���}��DCC�Bk<d��%��l��%�����Ν3y�W��� ��tf>{��,ʦj�D_��L���4}����-��S� ,i�P�K�PL�$�?v�J9� ����ƢM�Od�F4��DلI�=kOH6�R�E�DaM�Y��GT�c����S.����m%�Z�#,��N9���z�B��%�ہ�՞�'ˈU��T��TU�?�U���bQ�T@u�Ä8�EIL�+�w,d�R�5�7/����2�����	in܎�'NJ�噠}���:I����k�����.���*��~��~´"�WjV�שj��XX_;
{/��o>K���Z����%RA*�ۂ��׫z�g���u]Y�0�NǇ]������_ -�a��l��9|Gq���Ɋ��D�����
'�w���� 	�>#:Q�3`�CP�I��;a$j����ŷH�9?W;EZ��D�aE�*��*�n�������q�[��W��=Y/��~)q����P���x{�ӱ�2�U�D�o5�x~�ߎJ*�d�G4�J�	iizWx�W*B;Vh��FΥ��ql�t �������}�;-����H��9Li���p\�d��<�|#���֚f��X�]��b65���h1 m+e�1F�ё�м)� ��p������IKe����;S!b�Ǽ�P*\'��Q�2�H!�y��u�\�ßrt�
ᗚ���I��܉�m�^N��*�r�>/�>*�b��"o��� (l��h7T��!z��*z�/��T�����,"t�r��������>'�sCY�F�"�az���o��lF���}��+�+2��>?"p��M5bN�L/����'��ZA|��f ������!���q����͝1u�bUI&:599$]Y��|~��_�^?�_hgM(�G�ꦊ��q���d�s����'����χ!k1)��S��?s��?1���#��϶�%si��w������C��x��Mt�3�W�}���S���z���)T���蘪r����p=��N{��(�v�w:T�	�T���#�
qi�[|�����t7����W�s���0|%�oLD�AN�����\v�<�]�a�)������Nu���+`�oB��45�C��oڀB��/C�w�Tም@)b1 ��
����⧝�Z�hL�Ħ��)nJ�%�_�r[,1U%�2�T9T�cgU�	��jJ��|�ā�qJ
�s�T�"�&�	'jX#0�z���F���$�^u��"����,�=R=�g/B�����0��0 �e�*Qߋ>Þ��I�U�2�k8L�k�fstiD��}x�%U��rb9��𹗆V�@�8 `����ІV�1-�̈��<>=9��j1����@kj"��__��ȴ�\L�$b�F�c����k����no�r�P���6���$�?��|\1O�:��'���8_���,'�
j0$]�3F|D�""��BR.�7��lܛ#p��)$G�.NR3}����ӳ!y��<羠,9���_4〟&��g(J���!�oU'I�"G>���~CP��N�1EhJ4 �I~?+^u��X�r������N��Ir@p
"�K~����C�pT������������Rs��d��Q���%��Y+�zz��g:�zV����R���_\�	�ˍ�a[a����SQ��y_^@� �2G� O��:qv��f|8�<D����+x#�o�t���:(�<��.`D��k��y�[����S�P���˾�u�h`)���Fm����L���2nd��;SK������q�ԗ�d��a �`u/��/V���/u���oY��l�Buq�}�>QӉ:�K�R��-�9���(5`����'�cDK��Gt]	R� "xR�a�]F&i��T'���g�PY3X*Gm�f:��~� _ۧƝ�j�u�|��6��{�K��:=;߸~p8�	�6�+kao///���PB�]
��dBbf���P<��2�	��������;�z91w�o<�gq_j���(�C�0��?��,rB#��h�s|x6��Fɒ�֘�Q�S�M.h�L�°eW���8ex2���9�~�a*u��1��37#I%s�H�c;��|��O�1d�z�������y]Av�ļA[XQ�����F$���}E5,m����d�����XΜb�]S;��̶�5;�2��x�3���B��Z��V�z�~�sւ:��3�(v n8�k:v�u�B�������y]����]|hZ�K��%S����T���~h�f��.��&�v�@쏎B8C�>�H�j����O�c����ԓju<~y�"���x����~���%���y����-�M�ז���#��
�aCE���NE�MU�hHNI�a� R�ܐ�<Wi����I� �S�t��8��>8��*�rfk��<��%j�4��45���$�+)��T�9G_i���H�ؑzP%��DMI�0��a�����-��KӵQiE�_u&U	Uk��T�.O0L�6��iL	y�i�H�V���W}�>���R��~E�w��V�� n/m�z��WkB��N�Q����E\��I[t��ٿ�N�07�?���v����)���e�+�0X���gR7���ei&���Ɲal��&۵f�O���{�pw~���y��4~�D��	���������y>>>�ۣ�����Rg����zT[o2�ͼ��q�4�y��N��x��eFp�\���3D��5�5�t��:ͯ�|��K�lu�����^�7'��=W�Eu�-ӹ�~ϨI�n��2U��}'h�t�d	F�om|���+A�i�D��{&s��)\�ў�a#SQ�9N+�q#�k�W��H�N��2sQ�=W���B"���G
���.�C;W�,^��K<.I��ē�bK_Qǣ�6W�M[}�D^�S�MԪ�h�蚉W�U�}�t����)���I-�npCh)e��s���	㆞:_�ܠ���5{�(�{���ф���:�q2���<l�����m��G����y���qa���2�
�Ӌv�>����9t�
��rU؊;aY��:���w���2t6���P-�7�pf:f��L�sro>�������[o�e	�uz��M#.�d��!���|�I:�y�ꙁ���2�I�D�i��@;i��%f=`�t��@�}Wq��?����*yc������+��pX�Ӿ�h-�_��#`#�n��!��L�G4��u�A)X����&�J�O�MƸ���?\4O�ٙC�jOb�C-����Wf+�I���U\��F�u=4RBZ�*Ն��������{�(�_�x�Xh*��@P�Z@��8�տTg���q���J��[$$=g��s�il����ы�]D�H"Vص���)(�p�r��g&^�$4r:�C�g�R�SWI����L���a�]�8F?�Ixc�l��5uY��vtF�w�;b�
R��ɓ�h�ҋT�?j�7%|�1�/�G��ni��L��'߹�N_H·l�I$�O���aZ�ݧ@y�,_����˗��N���O�~�����/_$ͯ�=�-g_���U)yn�0��#b�@�j$~STTTh�S
_�vk���7%]6t�U.䡥�E�S]�?��ww����D��f'uہU��f�5�˅��a�b�����)g��nV�P��5����E��1�D
����xQ�G�LM�G�x>l��"d8ZQJc���R*�/�;���T�K�s�`��~)�e[�4G;�H��h�F�̘�sP�q����Ôz�VB���,@i��Ό�(������P�T�˺|o��oh0��MZ��
^��/M��5=��C���q��w���vI0���ri6�k�H���<\16��V�|:е=p�&lٟ.״H^o\N�^��x0�����1��Ù���ޗ�B^X��k� ^I�n��/[
�pD*�F���߱�4j1"���Wɔ ��U�1���
���Ɣgĕ�C$-�BC����� �5d�d$u��@ 4��B�:���\�G�-%j���]��ci�p1�R�qу1 m[�SC_џQ*���� ��^Fm/��v��!��*���rj;i� �S�ln��޾�Te�����nˡ�g�a���?{��3��P��pPBq�ɯ��	��AXF�z4r'Xc�]�3Zg��$�r=���a5���M���z�$ܗ�D�
�t��A/�:�
����ycM*����v�x��i���z8}�O�%C�׫�liZb���/��N8���K������`� ����o�ֵ���/{ci�:���\��5�u�8�n���g�����?]�C6�Z�w����&�*M>�D
���=�L���a��`(��M#Tc�����E�[Vr� )�@�"YE|S�`w��v\�]��ޠ9w��%X�M�I�9�Β�ςm_��{������s��.7M�*m������ۄb�1�v�@�T�����b���V��	f�����z��'�T�w�q�L@���pY����B��4sRy��IypgZ�s��i�w�&(&���霵����ÿ@�9	#��=	�p�q�̀�H�K��j��B{�������1ּ�Gy�)��g�p���2Oݷ�L3�J�������5�'[(2� �ğb��[@gW׽�.?�I��ק�z�ezc�R�ں:��LI/;���	nD��j����j�����~%�ؓ��Ģ�"Q��Uѯ��^��.T�l:46���!9oF������l[���#��Ǉh��~Q��z��T���A�_.�S��Z)*�w�q7~��1���I������iȧ2��zu~��ѯ)RˡvgO����?��rC.da>���KP#E���.h9-���d��_L��ɜW �U����z*¹t������:�������\SZ���(0/��!x<�������;��#O.���%�����5�Kݏ0C�PW��y�qx;J`q��a�������V�b�nզ����tb�Y{�9aO�V�����	��4��ja�J�^<��U�E�?}��4���EaɖЉ�O�[]��e,L���;IsN9>�l���]��׬X�,g�p���D����df_�A3H+:���$�{.9���a����W���>���.�K	��嬹�\�#B���8��r��P��$�����H�G���O�d%�P%D����-�N�U������_�K��
�_,��\;���д�~�۷�LQ�d"P)>�$ KNk{������.�����T-
x��������0xC�-Wo�:8O\F� W/��'T� FQ�H�:�viO��XXO@�Md��`��Da��`�Ŕd?�׉q��E�&����.9�q���3�����-�ѧ�Dj��C�j�@���1sq�_ox�E��s-���ѫ�yCp��O�7ύ�9[i�v�Pg�������!{���,Й�JLć�<�̕O��kЁ,��I_�l�㱽;(�XnA�~T�|�.��S���̴�^��?'�Lj�F��Fv����ʿ4C��vZp+é7��{�YKG��:YKP���h��%8A}�������sp^C����ƭ���Ḯ�c:�F�� �1��y ;A���2��hӼ*��*�Wb�WV���<���+� �x82<D@�Ld±�(���j!�<�Ӗt�d0j����8�B]rְ1�A���&��n"�N�q�DM.O`�v8�4z-�
�5P��B�+o�7�:5��I���.q���S*��aZ߬��K��q��:D~^����о�YY<�GN��̻�P�[��j���ލ�_H�ځ��*^�1Ĳ�w�kelw��������ߺ��H1�j�X�<ϸz���p�2���Q�EuN4-�<���ܧ'��{�%^�>��'���z/]�'mnV�������g3SS�8~n�@�	�ޗ䤤����v��Z��;+��tT�������ҒpR�]��bē17{"G�ӥ����U,��p/8���F�jR��,vN7�`xr+��FRW3BƱE��	O)���I��F@���,�ŕz��h������)�n��G��{�t��dc�i�ݷc)��@_�]�k�N�B�i)�T��o0�T�����e��?/|n;��c��J�C�r��*�8��A�y��S��O1V�f\���c(ݶXgM�n;�L�.Wlal��1��ri��Z�^L{
�"�E��ʓ��l�,����]fQ}�Sj��׎n!��K���~3����g�Z�_8g�8��m,�?�kbYXSf"������/èE��s�b����p�/i���Z�Q��Exnb	3#~*����}Ԣ(Qr^��W\}U���;`m݀>a���<���(!��K�H�yN�����u��^���R�Ux�8�P��8��n����Ob0����Q�~m����v4A~1ǭvS��υg(Q:�I�;'�d1����K��h����f�p)�=x��s��,3Z�l��Dѯ:��:��
����1xv�ĺ���Sㆇc�?zG�7�� ��"U��9�qn��X�O��F�*I\���آ�+S�Q�F5%���:>ъP�<�8".��Œ�(��JЫ�Z�%��i���gg�O(�k�8@�x~0�G�[�KZdD�7"��>���~�o᳡sss����\&D�Ű"��Z�G�A_�*�ڑכ���[wu2f�:��j�m{S�q4�{�Y�vXyb��Q4q��_��'}\1$4����O�d���$6���XA�^G&D<��D�r�\��S0d߀� XT����YDS�����;t�)��	������m��������Qv�V̂#C�e�Uw�_
le��Sr��"̨��Iߐڸ ����a� _t#JJ�97>���%B&í��tN��+�YC���TQ_�'���:X;F��ֽ|n�1j��Ϝ��Դ��ȴ�lg=a��Ȝ����~�m=�Ȳ�mN��9[i�<$����o��l��GB�vo�\"�b�j�T��Fߘ���FaP�Z�a�X�Ec�;6,m���M'��G�䚦EA6)��-!����&������@�%$}��xd\w�|z�v��aEy;,c�a�Zk����9��'��XTqg^TL��U�^�����R�� <��W�%��9�B͆R՟���Ҕҍ(�_r���<'�` �h�Np�7��4������E�d��*���2����z��8ǘw�����U�y4��[g"ޞ�uӼ�P�߿I�{��qF�+{�J�8vzۺ���o̻嶘�s�HʷP ����o�����òb>L
�L�e�~���Z<��-8�K�ڐ�Oѽ�l!�'(�2K�������Ѓ�g,�QK�j��'F��,)l<�0���1��=����5��CnX,���?��
��DP��������i���Mx%_B���`�����
r)w��'�}9%������-�B&����=�h�;�L�"���.ZJ,;�VQ����M?c,[l]\k)1/�q���'L��F跸� �[N��a�9R��R*��r[ZZ��u���"��z_,UnI�ѓ9%u�M�%d'D�#�3����{L�>���	9ѯ�o����&
	4�F*����c�
�i�B���/�Uq��A�!3�1�~�NH�\a*Z��7z``"֊V� c�`���
��MG�9|���-���`X�wV���m��ӟTEm�|\���	������Lu��Q�Yr��Иց-�ɨ��8ˋa�;�Q�W��,p`�w!G`��(o�+��uɴ`��9d�V֭�
�m'+�q2�������Q/�갋���\&<$(W1��~��
�{E���K鸦ͳ� ���[04�����(&t���Z�r([Yl�]��~�J-Ϫq�$�Ԅ��\9/6B�Ụ�]�>������vY�3�{��1a�m�q 4~�2 �A����d"���)�'5JJ���
��͜���앣T�� ��ɻV�恙a�� �i8}$��!p�j�UF�⻼2�:ϙ�o�Tp�ma� �a�;�@mN���܆QB6�n6�E ��E���Z��pL�5\��c���:O֠趔��V@�k{`�d�Bx�a�Y�jdk8+8qo�v<�K�����B����,��N���w�AA������I��0]7&�������	��C)��2-�{#~����{�ap�\6������1��(�܄%T�R��{Ј��,e�˴�x�d�`}��B����;Ǯњ?�C�O�wU��kBX]$�W�1��{���T+��d�Ř�jVlg�V�u������)�`̟t~#�Ɂ���*�l	Y���Yp�p�Q�0? �����	��^0�C,~��<P�����&��_x���UU|r���smy<S��io4��Dퟨ�Ɵ��А>
��ikk[�\��E���PG��/A(�����,屍�6bG���U�P�^Ma��0��S*)�	��Ԍ��?e��RCxrɕ ����Zb�"�}�*�A�W<<e��s�?i27S:��!u|�x4J5�G�A��r>	�3�BRX���m�)0\v�X�Z��qB����s��l��`˩+JZ�q$8��q��x�+	����4S�e¸a�uܺ�����@_k�n���:�I�R_����0��CNnll���4�7�UB�T�w����������/��:E���;ޣ%h�,��"Ü�j$�K,��}�S5)jt,��Ag�:a?^�"�D$DCЊ�4]P[]���N�X����JqwwNp+������݋[��.E���7�3<�a���{�컻g��1}�ЈBX�܎Lt�+goK�E㣋��:�4�2���0)&�ޱ8_������ ��3��zG`OJj��S���3~��T��dA�)�d#��%�7�mX�Ǐi��' ���,H���5��Y;�[�W���t�|�O���:���E>�_%U�o�<�#�N�ܞw�k�Xf�iAQD�I�Vz�g����Y��pz��~�i��w�9�d�؄m� {R)�Ze��3�s&��|����Q�Z�抸\����
�]#v��#M��<Q����.��;οaO�A rv�<��a��At_Gh���i������V0�����vHx"�o�swU=B�w�c��&������yƟ��/�!+=nO�M���a�S�����J��	��o���J�+<C4�soi�y�.zCCCO��U�R�/����Recә�-����?��;;�U�~�+H���,c���c�(��U���i�y�,�[
�Zh���W(�gƢʠY{�#Iʧ��;�3�Y���.�����~0:j���d�E㍺�rq�X���s�(��z��%L>��)H*�C#iz��!�q����})ؕ������x|�����v`���H������@Q��mr��体i.�^,,F�����c	��յnW;��E�2�ʒejK/�(9���s�V+E@X[� �����J���l%o,E�=#���_N���}�U��Z	~rB9-�}��tB��W���SV�axTtpQa�[�v�;*�Dݑ�c����'1�5sT���Ӛ���$.�y�y��L��?�xxxT<]t�RRRjԛ�1��0����P/;�P�ز��77m��teΛ����ل�\�����z�z?���p��J�~��Y�y��x���4����媗>�؋�U,vv��|y��G�w$
����%ilP܋��;��c2q�3�~'*J��2��Q�%طq�4���Y`�� �0�5-L��s ��Z�Y� �T����u��ʟ����x@B�y)j�G}S�pߏoLP�8���O���mن�@떡�=�tN�C�,�þ�f��\.lRVXԲ�
�z��O��vc{Rt��5P�N8f��� o�>!�������P>M��:���M|h�����P�IH8ڢ�ȉѧ���;NeD�U:�P;.\m�,Y�a)�Eˬ�U9�
�a"5�E�bD�B������M�q����~I��d܇�����Z�[@�7f�Y��[H<�ص����O	zD�t�L���6������g5�)�ݒyt�����[�l�	:������Tu����Ǚ���k����ϣ�3�f.m���r"*�>]fE�7�d*o%�Yx��c�Cb�����(�D�U�8��X�!���l��!���Np��{ؕ?��0��N�]˘(�Q��ڜjo"��.b,�
����2/e���'^�ځ6�>]|��F�ʩOy�㺜�O�mv��%p�.nD�s�eh���G���8Mr��W�4�@���:>��'
�g"s>�G��㤿���g:;�X���v=T��RyVso"������++�ǾųN�,,q9&��s���_*?��QIߎ���tlg��������5֟WG%׌����Z��h�=�f�6����k�g���/����\�Z����[�4R6��Vm\��y���uܓbԨ���1���,&�ڊ������;)!��+�ظr�o�l�*c�)ރ�NS��3��'=�_�(�����I�q��u����2P�|"��1E{�@���FOwg�����|/	�5�>ڛkBw�ꗿ/^��E��7�b�7���?��:�B�����R������3|i��VJY^Br8�w�C�ۢj�i+%��_"F�����cc�+{*�9[xf"��JR�¯晘�?�ޙ��!��)�'�}�� l�:+;���q�����c'��%���5)禜��6���Sl}e%�2���L��H|vRP�g�@Lh��Y�̀���Wو�6�u�a���;z�lhS��uu���^�(�(6�-X~k��D��1^���#7��UaS���O�+���������T>B;��5>k)�Io}��]�bC��#�$7ps�^�\�;�k-+C&��?T��2�`����Ӝۊh�����t�om�9��:&���F�o	c2����)L[Ƥ$�E~m	u�*��'���)Ym���(��T����6�?ړ�ՑB+ۜ-w&m9.{5j��_Fv��w#��O�&,�Փ0��#���]�n�#@{z��b��\�lkû�/��H�,��o�C��BTupå%��NF�G4���)%��Y��`��Ji�
^���Z��	�	��#6�����6E`[�d��P"���9-��_��%2���0,Կ݄��^Ƚ�f����X����k�6�~�lj�,���ٯ�4P̵�=GC{\�6��J3�x߷��;��ݗ��e�.4�������D�lI�5�1�����=&��h<�]��IF��YDCaq�st�?���a�k2Y�Z�������멫�O�y�a�����>����>�u�Q����G���.Vj����~N�'���F�6=��!����ULD��������Z�\���R�j���=��ЮҶ�Ʉ�L�>�����<D��޾|�Õ�c�Z)ܚ�7��G��ŀ����r�fӬw���5�И�]����� Zl���>��݁���������y��1Ru
G�_�01L����k��1Np��W\"τ��a�T?ey\Q�ӕz�Ơ9��'Mge0yM����D��0�<�_{M��@f��V�vh*�	�Q#��'F�.bHtd~�k���$ä�ץz����rqj�;1��7D<����ߨ�,bd����'#��J�o,�m{4�d
g}�_I�H`���/�my�[s8*L�o|9�hw�������mG@��� 3N,����(�y�Q)�כ�v4c�g��%}��F� �S��ĥ㾗xxr�o���N��7s�|�p��#�#��-zh;��g|hub���¢bV�͎8����9ih�#���qX���|�Ǻ	�$�����P�ǽ��� !܎-]!����u���{�!�Oc�3nwن�ҷ���MN���������~0���t7�X������m�eґS��o��=̹�������G���%�Z�QV��u���2�w7\�L;d^��x?/g�Z�?.Vh����;h�K�L
 ތ��)�X�h�.d!(�U�7����e����V�K�=Le��	�݁��C?�І�VԼ��������>ww�[N�q`>�\k�zm0ⓓ�"��A�����~cq�L����#Q�k��L1G�bB].�r��B�j�e
������ tX/=�>\�ԙHn�{$�m�2D��Xj�X}��{ڟL�:�����uu�7�cZ�::?"0���b�m{�ɔ��F7��n����Ѹ��Y�ƦEX���f)���(s���6��y�,�j��h��[M������i
ѪI�����D
POf�i$+��E��$B���e�C�}���z�\��h������}����E�D{ME�Q.D������~M���4)>�g����B2b������ {�;e�#�d�\j���九�zՇ¬�Yk�=w���g
P��o�m�����T������-L� ����,#Cn<l�� �]Ո���-7�=�[�~]���x��R�@rx�Q?"�����/�m��T�^'�Ќ�E�5.O�&b�eX��W�;:ΰEpm���S��[>C�]�3�P�{�u�rO8��9� pY?v��\��],D;�Փ� TR���E��������r=r�\����J� .o[O��=��Q�zQ_O�vs�\�)�ﭳ��c��fc��ts�Ծ�ab�2�h����r��U�����q�ԃ��_zt~8s�+��vRUn��3\�n�-崡�bF�\mj\#0F/��N��N�-W��AOg>�먬�r��Κ������0�V���9$ٵ8��¨��I4�b�lDN�;�s2��E�'��������~�o�h���*������4����9����ׄ�}�G�	���薕+9�=�BƔ"��Ⱦi�E[Y�mˠ|	�)KI�V�#j��1�e�Q�;s���`���@.�A!���:�M�7��˳�*���������]5����O�*x'�f��f���-^�����yff��A�k�@T��̌�]��
�������FG�>�o�F�-��^�����Jn޾�� �pf��I���NE��{I�?�c�c䜮b�0��p� h��Ą��  ��x��n����C;"��ߵv)@�蚥 ��#�M���OF������ ��/� �6���?��\2����p�v6��&\Q�s�3b8���3S�O��-/́�c�*�	��j��������9>3Z�K�M�u���~�7�	j�ŝd)1���� X�ЩJ훓��j�[�fޫ��K��x �k��E^t3�F���C-�^��L��q��	�'<�=�|zM�"�%W#�1	.6C�~&0W��"�V���aO�\x,���½��	�,L�I�E��Ӻ)>��1��%q,Dx�Q�w՟@<w,�|G�Z��l)�0Z��Q�%��gX?��X<Y�3r�
8�H80� Vʙ9�1N�Uc�U�4�H���Z���r�j�G������$�9��YW�a�l�ӂfs�>�\-��\���-8�A�.P�����ؼqد����������)2Dj�B�$5R�޹���v\I44�Q�TCg-_�jt�x���e@��������� vNti�f�G��5&p�d�C�dl+1�zUB�����=�@��O�����T��Gqx\�:����� ��+j�;�v�Z��o�X7��3?|Zϖ�T��ph���<�p��p�Pn��G�>��(�h��,��J!�͒�3��{oB��sJ�_��}���l4g�Ξ�!='86.jx\�� ���zM8���������D����Q���a� V	���gXB��M�Ĥ�uZce 4�?����1��bJHH��r�}���u����4��X�7G�n>�Y.�(��[D���M�������yI�~��P��ZW��0���Ѽ���<B��Ub�W��$���yj�ĕb@�C�	Ë�NB��}�~�-�u�;�C�rc�v`$j}M� �l�q}�ςI ��kw��
��B�u�@�!�K��{�]�K,��4D�#s�N�:#h�JlU���'�- �>�Vi�=R�n��~����GBlw�9�{�~z�1����4�Qz+Zkd�����bZ����ԭ�­4�x64�7ƺⶥY��/�!�Sճ:2�6/b��zډ���O����)T��w[4����%� ��!��~��}(�zr�S���B�$k�z�Ju@x2V���â�7@�Ӵ�'���yxx���Ճ��^86=/:�&k�!�3���-������kn����0BI��N��/��̮�5��K����̚d�#ʁG�%��^lP��︯��۬ث��~�q�˚�Y����O�[����l�p�:��������_QY���ļ�1��(���]�B�Z�%�i��o��@��~e?%3�ј�]xVb[�o\`ڡ�/�}��ήC�{�!Ϝ�ZڱT����Q?5u�3(l�]ɸ���=��[
�bO�M�û<�n�#��|w]�a#���D�%�5'A�kv����'5ޤŖ΀d�G����X�&j8����6S+a�?K�:��;��0s�^.jM5s#�C��{�_T;Ji*�m�4+��Kc����z�Lrw@rF�Ȳ����IY���N�����r[&�?u4�&>6����Nx��0�ɭ�O�$&��e�m�(�BϚ*�h��V��=ծ�
rI��K��2��������Z �X�O-~}7&:c��7�@����CPF�X���lI��H��2�(��ð]�?f�@��yVik_���71�<��Eë";���߶c�@	�E�$��uk��T.��߲�Y��ӂ�6����[�\� ?����}4nt}XQ�*�pIF�u�X*Φ4�q���ډX�㞿.ZCT`��:W�*>�vUO���뚈�Z_��3��mOJ����a�Dw�î��t֤�A�0t���C�r���sK�qa�1�Q���{���o��й]�`�(�tv�9*��]KC �_40bl �1�߾ZqH9���u)��{�����3f[/?����1h��Ǿ���Gq5��������*�lT����4���F��yD�(���<��S.q��O������\8f;��O>���U%m���BH�*&:)�%]�lH���Wi��vȰAPX-c/
۞�`�T���B�A?�V�ә����|i �Z,AG�X�88�B�bH}��iv�}Qn�Ҭ����"�K��s�v��5�'E����R#�Ƶ���Vy� �*+i����̓w�p\Z���x@cr:/���@AM%Y0wQ py���I���G��m�S���o�ڂ���k+b���1�S�A�����9P�A�/�������a���B�ŧ,�)�iJ��SR����`u23'�2I3v����,v.��Wy=�8F5�ص��	ۢ�y��(���>$f�ASIЂuҪWX��л \������bM��akR���m���n�A�Q�D�j��ueMj�MKt �j]\�Y��;�Nrt]�6�տ�{��HO@/�\��_��o�����nO/��@ �M�@=h2o�\��M5b	��B���ͫ�����o9�{U��2܅dU�Y�RƲ�Ñg���$�Y� �����5�_�.�� �Y3��7<��%�8)׋��U�Nb��ʭ�Z�Gp	M�_��s��~**Ρ^���LOM�4�����Hu�a:is�KDq9���=>��8)�ݬ6��
)��6I,0�q8u:�8�� ��G��x�R��BW�=�� �1���i�36�cX&�Rh[���͈��`Dk�� �&b#�+��D��Da�l2F��(Q��ȇ�]g�V%����o{1a��}��C�}1�<VwP�2/����d�35�+V��~����P#T�����9a�m�&��t�� �F���IAP���8�맚+đ�|�'�W�w��{�^7���wi��N�I�aV�1�BD�j�3��E�N�q���-]�BIT�Q����jd��- �o
�>����wM��dce�4�\8Z���96A�1�78�̹��ᨊnC�Y,'C�&���w�`+l{}L�P����S��x�B��ڵi�K15�^3M�&`�9��^�0蓬3h`q@;����g���>�"\B��o�ܹ�}����Ȁ[���'���۝��+��ur���*�����[PG�	����7�L����-`���� ��CR���7)K�v׋��t��ק����h)KFQ�X���T�L>���>݆��\��qQ'�U,^��^��*�I��[xx�!A�茬���F�(�����(�����'�O�|j��Q�����T���yv�௡�����CqY�y�q�7BJ؉S��������މe�-��1�~����fRQ��O ��C��s^�L�W�U_�q"�s4��0��%���2x��7�i+��F-� };s{�|#���(=8~��$�����.��.~��1����bw Tq���x�C��"�,���z��5�'QLT�֓�v�,����$�Z�F�dםi����Ƙ�P�#�VQQ8M�����"��%�5�@����z,�):	��'HrP+r������w�mpK�r*Ms"#��
VSF�ێQ��/�#&�6-�~ѡ��?��;��g��~���l)�w�	i�}Fv�K�A ���۸��d*�c�IH�w��'���t�w��M�CM�D�;��>��>��:��!3�!��Q���c2L5'RX A��/��G/T�(F�m���("�A���Ҿ_f$��ƓiL�ņ�*a��1����O0��0$$�OT��_f�I�؉�ᓪC�j�7zbWp��6Bql2���tZ�Z�8��vG�N8��kR���#&�MN�I��R�c0�`#b�}����	DIY�QE6)���G�JH-���:R�!`�%1�=��ի��a��<���s4�l[Λ��M�ǃE�o��S?����˯h���`��f9��BKK۳]���GP7�����.��!��.�QeUU�]O续Y���M:��i�=0�ĩ�1$LH��bJ�%�6mN�υL[9X�d܊{3�%U �^)�o�ff��s�E�Jr$�Qr�y&!H2�9���r#�:6<�Ut'J!GǨS-4k�{��e��� ��>Y[&�C��غ>��D�����s2��S��?���k�����{����2�t{6\aU�6 T��f������|���\H�	�������˰ƍ�%�����ڼ���ͼF�,|�|�2�YlX;dPv�ǽ䎻U�R�|���A��؉^e�f�"K��?��\�r�71[���JJ�5��kS���2)ˉ4�v3�M�m�Қ~�=~W:8Y��W:�u�YE��G�A��<ġ�?�z:4Vm�5�a�7��>�(6�D053�h�?���>|f��� l"��!I���g!!���tdI�W���Wu��z�-$�Rnv��o�� �ɹ$�_}�<��9�Kg��'1��6#�wK� ��#g���/_���pkxg��
�w�/�~�{_mu�@I��D�;�̦2�@�U9����?>��T�+�C�Fq�]���D�r�zgog�����A����[���?V��k3���w�MX4~]�M�%�o�>�	N��f�<���!fQ;���M�o��)����Y��`���6vO㧈ڀ��o�=ή���}�.%G ��(U��6�6m�K� �:t�5Ej�k��Ҽ"��ނv��b��ro��Ǜy��s.>�j�j5t�o�'RX�?���7#��H���Ug���r�Ў��:�R�咮�0�j~- �g��=f�ܖ��u���i��0���B鲯X��[��e_1A2�$����I����r����T+++n�$��9e�w �$SEUՠ����о>QF�k��P,J�, �ʊ��(��=Q���kPo�m1�7��N�x�0^���q�iܷ^��}o�+�Jxt�)��)��</^#�E�C���-�
��j��͵�,�O<l5_��G��
A2�4	����6��&&�	�
�̏�#�)rZk�U�Ց@&�'���-k�00��u6	�'~H;�ba?��;��������RІcE��J����eNQLɶx��o.���zۤҤ�үJ�_s7�CQ|*��z"�r��8�E1��ZcH x��	=��ꎗ�����PP�O�� ���-��]|�{%^����vf{c���u��]��J�6"7�]�5�x��ĺ �5��!��{O�e����ʼsWNc����!�" �����	��Ɯ�SDPWu���w�EP�uT2#����s���$\L���n$Gm��֎CY�)������8^�z�>�BW3B���S�# H!�쵇�Uӂ�*�hB�Ā�j�U�9m谹�;b��4f��+�;����7J}�L����	���KE��y�x*�8��^"&���i���H_���R�v��pRh�X 7B�G1i1��������.��M�"�|����
�P�ň�7�6\�>w��B�(�X���z��7A5��VgO��ى^Z0ς�����e8-	�fX��>y@I~a�ݘ![�)��i
���*�=�����R����RBmi�kR��Cl�EP�$�p����8�J]A��EV�J�QC\�i.��jh�.?C��k��P����㢐/LnC�����Lg�� �� ]���4$IbX���g��˹<@)Ma�����$�e\�s�Y�M-LcU�h�A&������cɸ�"�@k�Jѿ"��C������~4���"�l95��"_Gi��J=M�����-�����>
}��wx��)��ꝓn���$ۨ�u
��G�ƶ���=&��w�U6:,Z��ŧ�R�G�����˲�i�cq�D�& �_<uf���r�g7����Q��4T+�P�L9���y{YZ4ὼwZR��6�M�oYڸ�H�����*?\�����j9�[S���E�B]���2V�)�!�2�wx��m�q5�o����\���j�Bw���ЙJ9摤^T��޺Mk��}/��$���RYh�A͙����r����#�r�:��@u�3<�K�mr��	��<�뛛x��*��8�d̐�u����ߕA�)�%j1��<�k��k_�=�y�|���q��^RRUm�]�[A�[���$��(��� �B��g�~�z�Lw?Q�.{]+`h�E{�n��H����ݓR�c3X�n��N;u�Ї�*��M��?O�acW'�e]���{��P!�{��e��]��Ô#֊�� �W�WS���v��2
����{�<U�����`���w���*��Z:	
`�fM+�s�y�\�0]eB��$���ky5S8�M"E�m[	��"���r�5�3��*�?{{q��o�|H���/���Y�YΏ��p� ��Uut0� �J���-���0h��L!�G�};H��m��)ۓw��yU�|�>Zy�A��-��f��I!����8�]������b2�`��
T�/��ϡ��Z@r��1���Wb���k�R�I�8S�(ns�������
����!L���k
��<�ÙZE_�Zxg�� ��[�(\
��cӰ�H��G�H����n:50}0�U���mRmT�*�oN�
��4�h/�����o�O���j6G���Yu7L�D�:�y@{�/O��Y�t-�+��X�=4��[�X٩z���ݐ����˟c���3��:�BN*�ئ���N��4c�1�\4��K�$�7u�gټ����b�5�K�)�n�l�&Ҕ��'��1?�$�1���0�̧�����0�WُP�����:-�鈸��Kiu���&�&���s���B�|\��h��i����
aRa"rj�+�,�h��x<o�PH�{_~����aҾ�����\��D�!�@ŰER�w/����?��y�t=.�zT�-���3��>��_��7�I߫��<#��U����`2��&��ȸD���v�*�L>�2\�QD�t�e�,�Ⲗ^2o�ZW��^���A5'��4���Go��;�����m�b=3�� �*s~��¹�����c;`ж�qʗ�F_M�+��}�z�G�6=�,��1�(�ee���A��_u�hV��U�t�%5J�T��5�|YĜ6�#�Z)W�󘘥x�� �!D�R���)g��j� 9�%W��7�~m ]-7�JWG�4t<��m&wD�ҹd�F�uP����&z6�����`�_�� ��	�l��w珖����(jv�]�Eԫd\j=�����]n`y�5�XB�%��F/�)�|2����������K��}<�ξm%�ul}��~�U��7�TLD�{ߢ3I�j׷X��5#'�ͮM�}v�S�M�
ٍcDd�4w���ˮ������Q��Ff�� ��i���( �H=+[�!��BS�Ͻ�D�MO�֏�U�tAl�!(�
�?�!�	G�#�R�
����%=�!ue}�nZ�=G���c�'ס�}��fѧ:�a�(��g�8���c������S��Vm�
�����:ߣ���9=��!��ͥ3�"8�|�\L+�(XԙL��ť�khD�v���^�1K ��9$f��5� �����;���d���׎Г3H.:	��.9�>�*��+Wg�$��#��GKդ���1�bTee}��N+?E�M��ܹ���e�(`:��D���8�d�`�����	l������Y'�ټ�MF&a>v��l5LU��I�v��m��<i�&��ǔ�߇�l�VǾ�R�Bi��Y^�;����,C"V�f,��Pig3����H(1�&���*���"K���U������G<Zg�U4+W�Gy�3z��|�2h�q���L��W��ׇɦ�a>"�����&d�,��w��aY��M�/�^tِ��\���YMÐ�ÉC�1)^�le}R��f�������4gU�Ԯ��_¡R����d|g�u&�Ŗ6����V�a��R.��&&bw���NS�>�|�곯 ;5�2�?.K�����+/��E�S4��b�ףc�����0�b(����^5��ۈ��$�fk�^��@�\e��@H���\���,���m�0�v³� �u�s/�s��������ݘ6T|���^GF}��ㆥt)^V6OCm��M;�A�?�h������|�B��@�u������P�w9��*oU��x���c<�ۏ�"[�JM�ļ|�LEٲ�DC��c�C�&|*	q�z��`4�����-��@r����}�R��ūaҭ�t.��v_Pㅺ�J��BY�-
��������R�3���Q����H 0i���8{zx��w"O<j�t����\�IN��RC�_�������ݴ7+�~�{M>Q�MMb]��]u����P@3x)���$�{5r���q����Xj��:7�Wm�����-&eN$p}��T�W��nT�?Q���`#�����/?�1��U�|��G�ؕ�>Y�V��Ņj^�ΐ�X'��%$�a��^���!Vr���ш(hi�cb� T���a���O�2 ��u�}�l:k#�pk*HI������� �Os���)F��S��4���&���پ��xL;�1�F���1�x�R.����4q��|��Q�d�i�3�$��벑���_7!���Tɠ
�z����TuQ�2?�92���\l��9�ֶu/��Ϸ}�B\eT���iM��Q*`4�*~6S?f�.��,�^E7���mP�*_e����Ga;�� D>GçĉO�[����n���jQȆ���<${�JJ���	��;�����G9��t��Zg�����$��^�d����V1 �b��xp�v�!�;�)���C�ph�v�λ�|Ԫ�&H�z ;eu��41q�Q�#+n�1��MeB-)���yx�}�+�$4s}��)�7��y��9��X�X���BJa���X�HZ#ԁ��J�O�)^��[F�XՈ+�e�R�ՂA�\�-B`q�e0& Τݢ=!U�F@�F�$�-�ڪU�ב���d����z�7����c��b����#�d�hަo��������{l�I���������� C5��F𡔄�����N�A^���y�g퐎$��Q�*�t!)�;U?��r�>����8P�z]��^�,^�p�B ���\ݐ�_8�O�׽7%��˙���F'/��(���[�$��
cO�]!��z�M�G�S~�K�`�����1��k���uQm���S�\33y�fS��b�vR�{���U�>�X�v������Z:$��3�Ijh�.����P�J�ʽ`�E!�Q�)�����]���?�&�}��n=*J�r#��Zp�K��L�{�H3���F%���qgj�܍����|�aK9���Mv�f���	~1g�zߴ��؎l
� �c4����N�#�W:�"��+#BX�}����J���o
������u6|��tKM�0�qbeC�	�J��ĥ8OP�n=,��lR7�U�"�vA�!l��Ye�7G'l:V�%�?d:)~X;�	��~){��B�Y����p��|�9T��r�^��Q�Y�N�ڣ�W_�(�F�]G/�9��؏(��̷ֳ��IsZ�F4`���)|`�Ԁd���&�e����Ƭ,
f�j9�Ύ�ˈ�2ۛ�q�q6���:�X���b�	BBB���@� �<�$S�5Ps���^\\<��+�t��N;$�9B�S贺�)��@Ic�5f�T��F<|�CȦ&�G�#��5z�7��υ��q�{����W��C Ω�f&��PS���Z�J!.�*u1<F�p����|/^^0�����bXt�|���O���"[���˾b�6(ɤsE�g���:y�����zIIK�����F�������WU]�mB�㖮k�!o]ݙ4��}s�fW�GL.�:�LN:fod�<\�Xv�t�q�ܟ�}	��X�����GJ��S�@��a{ԁ���^0����ĭN����:����Wf(ʳu��ه���};x�b�o������dM���V���R��~eQB�|v�"7w|o�_�o�`Uգ��2�*�n�̝����rQO�Pq�-���Sss�)�����,n����*�C �V�}��#٧~�c�C��+m�75��c��\�Um�����~�AW�3Uo��j��b�>�g3�x�D���;���^���NG��\x�P��5��b=IB��b�����#$�����h�E=#����r@�汋�����W���~"\���Y�7þ@$���W�r-2����%������O�E�_t��m��x��<f��͔��ֹ��dY�NQD�JN>�1��Y�B�����6�֟M�$�=jT��r�sd��AE��rz�zg�`�w��E|��rQ�B��➏||?L���O�C~	�krS_���z�}�2t���C�?��9hX�x�[����ozV�ZG�[<
m�t\���^�@Lm8_$[�.�8�x����������/�̰�8(F �*�:Qѕ����w�\0�j!�HGjTMP�5�9kU˕L��7��Y�UB�臉�d �k��<e����� e���̍�0e�J�:δ�IY����� nC�(�zC蹧�~s*���Z,�
̓R9�����VTDj۶uz�s�Z�C^����5bI�3
7�t]��T���w�	.$;���G7:�$��NTf~{h�8����������4E	�` ��H�c��^��t �Eft� ��4~w6(`+$&�\����k��K�EL@�������ۛ��ˍ1qq�g��B��i�u*�8 ���\��}�۷�9�~Ճ�H��::���N=�=/{���p��3>J7���d�r����hw(
��ZZ��G�@%�O�S.b�Y�i�֭}�$�-WCD+��ߤv1��ƻ�֣�m�|�T��v4���->�<c"���	�Θ��U4�Ta�S��`M��`�9��(䁘 ���(D,n!��> �)S�nR�gEZJ�|&��p��=Yb����nj���������sh�ȁЛ{�R������!9s�Eu�abbb�^�a?<��D���x$�N[
f��{��ykHYYY�s�����An�My���p~%L�0�\�'s	s��t5�z�x/u���0�}~` ���k<	:ۙ�1��\4��p��=�F���|�����y-���諸_=+4q�ЉG��; i�pMV�!��5��`�Le�|��~{ꦎ?s��|����z����`���(TbL$�
��s�c�|�X"��̀a����J!�e!���nT�NMM9�JI�v0�;l�*�_�N 23��'i^ׯ�~a�f�y�j|�N�
�y�䣬ʐ��^1�j(��;8 ���!���ݙ���p�~w�n;�y�םF''A�ӂO��Ff�� ;55<�u��֢1�.
���b�t�K���k���3���$�ͫBN-��S2�)����,25L6@�:X �\�9�Ez)$�N�݃�ccW("*Dm ��^j���TO��H��ч_�vPA�M��I��ڌ���A��z�P�9��^�3���xT��;����=BAA��������\$�>d������d�fi֛5�ԙ�R�7,� 6]dյ���^�;6+j�B���R�|�2j[�T?�1ax+��(�\+��~�8�5���ժ�ުYr�$y�?t *!%�+9_	CUˏ��I
::�
�{��q����,b��4ޞ�~;s�Q����)�Q�������|ZŴ�-q�z��W���W�Hl����t��2 �<�o���`/Y������ ���/��b���4-���))	���4�X�)/��S7�_)R���Cb�F�9b��4#�u�B&1����IG��'�S:��	: �0�k���*�m��e���ᾟ
q������׷)r����ƛ����p*��qG�4,5��U����(����?��' tc�����6.�I��Y����B�m�5�M�(*b�98�/U��?������`��Hi?o��/��=0/����Q��St���j�Ge�m�R����P��򧚱�Ώg֗W�`2S�\�z�
����������|���@~��G��'��~��R��wH3B+��;��ʾZ*����~9�c����s�P����g���.'DZ5�t�d�naa��H��h*�W&�-��B|���|�����Ŗ�)��C��˅�4t]Z��Ў�-M��k��۽����Ǩ$9H"��cQJ��~�;����x���zk�&u��U�}:�zû���}c����������b�4H�_^ ��Ǝ��og��/,0�)�H��{�����I_tӎ/����NJREh�c	l�|rŰ��"�B?��K��v�.�@�ot�D�h�eee��T}TU]�6
��HwwJJ7"�Hw�t�t�t�tJKwwwK׿�������z���Z뉹��h�v܎� �wH��{O0?�L�!J����z�!�HR�gl�T�&jZ�_�#���@y2�l����o�tc\@�ظʉ6���=���17>�K����,�|���1R4~�;���:6#C�UX�*jj<ey,���<
�W��J9�5o�b�'��0L@�%,g��Ȋ��	`�����w�Q��;x(k��s�O����u�J��P"=XW�>��_��T��u��L �|JWsլ�:�:�b�����D�����̖<�n)���,R��ۭ��C���4@.&����ϯ�'gs�[����m��&n���z�dh9f�`@!g�ghW�k��^�a
�T�>��i4���+��HZ?X<�h�ѻs�X�� � �&m?)R�ٸ+��R��'�����! �&}��z�5��ji3u`���a2J�������P��KDЄC���(l���r�}x�p��\ ���goA ^;��!	̩����!�� �D�A���SW*jj��Z����W�����zt��!a�ӿ����}�f[�����nHK�q��]:^iD*]-��Q��"����t�<����\B���WGr��T��)�k�ZO�~X���,��u�L�^h�y�b��Y��M��A"�uTՍ\��<!AD0a,�a�����:0wG���߈W�ښa/Ӄ��������T���#O��Y��D�N�+����y͸;¹���fE����1h��=���������"k��s������&���f � ��?B��˾����h��q���/ǌ��[D�s#����i���4AN�����^�K2��p[46V������->(� �?7��,�����X�}<��G�r���Oܞ;#��1h�J���W@�F-�t-��@lvs̆g��Ԯ|�)�{@��O�L�v0�:Jw�����Ą�I'��Q�F	��ں��,������?�ׅ�3��[-�'���f`m�ѽM+U*Y����ݤ$e/�DmXXx�
,����!y��S�����M�C�ɣ*(���!h�����w�ih}��� *��b�3`����yы�TA ��.�(�l!�$4��O�v��ղ�|A�?`JZ�6������$tئ�&�c�өK�O��v���rS����E!����������F�gNz����Lϐ [��e��'�,Xf�s�%��4�����Q�%Ψ��dfʥ��e@��R,jQ]���!i��!}����&K`"!x�)��xhhh`` ����olW_p�V��]�(�l|kAJ��J����=�r�����/��-ߦ�~Yĝ$�mEr^*���9Z��ȷ��w������]�'\��z�|�\�q'���`��@q�� @:�v[_�Z�Fy�~�� 0��x���CN��o�h��0��/_�Ė������!0��(�l��/n�^�ކI�����5dl�m�~�TQyH��n� �q����Tt�fXKII)��� 1%e ���/�aC�T�p�`��`���N�o9r��2�'�ù|��u��|����7~B�M=��;�:f�������{�#8,:=�Ƞ&��|�mP�U�9����|#�����K��xtU��g�G&�f�ߎ��8��֙�]��&+�[��-�MFRU53�;'/�2��)�48(b:�բ(�qFGw��� ���}��R��bm(0��|���i?��R	���B��<�o08<����6�������x6L5FъJ8ݮ� f5;����ܠ?�Xe�(�<c;�a8�ww>�i�~wG[�څĹ<~�1a�`��j̴;I�����S_4���7�� ��V�v8�qX��H���v�R����ܫ�?��g�s��A���м(5��r���o�Ǜ���w`��"k�4��uݖ˶eE�� �����/1@�y����G�zn �r��	v��|�lGgU�\?�8R�#��Y����鴥�Y�]nEn^ݧ�f��8��f�w1[/s��y�]�2{�L)��6t�ϹO�����AC��0�(����\�jH��X5�h�8r��f(}�x��`�Ւ���ƀ����r�j�L��*�u۵���m���o�(�
���xj	����EmٲEΛ,/hg�pj��?1�K��׳�b���C^�ӥ��`��
<��\0P��=8�/��ol�<]lh�\�[Lq9���y����"�{�z�Iږ#O
�&̀C3Ԙk� ��=v�#�wp8Xiq��G�)Kg��ӤS�����X�������;�G#�0}��J"T�����1j|}y��<=�y��s�M�s{8(�	w��(�͑���������l��@.M�[�?k�^Ֆ��N!t.��%o�{��O�/�6���_�ò���2����3���5m,������F�_���1Ŗ�b,u�pS�}��������I�����ũ�o��tɝ=I[F��cJ49�M³n����}�G­Xi�P��ٴ�^Tv��
�^���b���q�������c�g��lS�����{`Zc�}R�f��]�=X!m�vբG�˒*Γ�/�87Q�����tGz��-ب5����K�3�WQ�@��������AN������
/@+QG��F37~���!u���ƥ�V�v��z�bh=�r������������?�/����_�����i�ܽ	>��m�W�ۇ�����^�����qɤ]<d7�N�N�{EC�����I�?< �9	p_�Аʯm�H�䀍�1����mJA��+@7�zJ<�0W�� l�]���24	/���-����Ik�O���D���C��͉���`�vd���ƈ��M@B[]s�El����w��ڶZԏ����c 2�n��L���������J���z$��M�~��f@����R0��ە�3 %��~x
�HC#5�.A�Җq}1�`���@KK[\Vqt'�'5���$m�3���[���&F��=�����S?��'�VJG��(��(��p��Z<c돒B�;}��.6Yhd|�)p��v�;�n�������e�1�"��M��&J��|AcA=�C$����T9�lY�����n|RR!S�,��^k�^�:g�-xV��Q�~�c�㧡�B�5���E� w�aJ��b�>��Rbq!�g��;�56_mx p�̖��b���>�h��BґY�ʐ	��T�T`�ɁRi5`c�U�|�k�HJJ���f�>�� ��*�I��y��ḿ�cR�g�{H���T�[��Q����yv�#B����M�O��k۔΀�ޜ��x$n/`64���&ep.�~��)T����H2����6���\�-o�	Ъ��ME�S?%�M0N����l\N�?䫴�6�o6�|�?x�זO(�����l�-�� �I��k
Hy�uPo���)��r�JE��Id�s�?WI8'�ˇ�Cs�� ���}�?A�>*�շ��=���0�
���\���60�9mt&w1���?�8%~H<��sdخ�2S�h����i���}��Rd�3� �jP4��&�����҈N�9�0� ە��[hk�o���P,C�
�j9fl\��q�Ô�R��U���2�����\b�zޡ�~ zJ,��w��]�&��4�?7�7���e,s��T��~i���h��0�c]�v�LF]f��G��[^}�sp�AV������̅8�h/��p��*�o00X#�@��_b-�''�u�X��irأ��&�@��o����;c�fŁ�0Xr>�I�>>�<��$�����W��P��1O�CF�_�V�4�mi��Z�N'�Ve?~{KA���yP1�[��,R�3�V��Ȏ,F��!4��s�bk:�2_�m��V�;�Na��w�Q.���2�)��'����=�dr����u��C�]R-F��6A��74�Y��KK%Wn߇����@��������`����=�}��|WZ�L ���0G�e������-�^w�Ϭ\ٻlw�4k�����0�=��bV�lc�z��l���.����,� v��/�
�:�=�=���'"��}Ԃ����:�A�C��z>���W$C�g���9"���!�5m��;���y<X�D���+��F�nW��s΀���Md�ц�Q���BF4�aJ�J*j���.���c|W��.�P�/�*�,�� 7��V�p=�@��J�𦥤�7��LO���V�)���S��A0���!S��V��延��+(~����8�I���	"�JLH ;C@pX/'��'@���Z Ӡ��zMq��j�������ѿ/��|�o����k�mK@(����x���Qma�t�Y�� �զ�8��t��� E���HN���I�ʻ��M쎻w���*'�3 4�ğ����"S�۾#�?�8�����u�O~Q�E`zY(ނ!a4	|�3���^�hM`�]R�+���i8���N��=�<�Q��噎eJFv�¬�����%��O��M%��ջgB�MY{ �r�m�U�k�Qr4�5.e��G�v�i��ÍJxJݐ�и��`Mk3�����pJ*��lt�v���w��p�-�U�#��rM	33j����ˮ��@���ZC��f�B;��1gPA(
i�g�u��LFv�S@tπ{=:�����x�K�6铓J���&���<$`覀�������'C�f(�ҵ�&��L��B�yB�����8܀���:/Y�����{�("R�-@g|�1���I2���kS{H͠��.��rH��ɱ䢧�O������tp��<3��a�U���s�2Ə�~5|rACfV��	��5�fW�u��%0יT�v�4~<*՟HyS����a�R��E��Z�w����ԼL���,od%���
��p{��D��'�(Z35�ww�#�t��Op��Ŭ=�����=��������;������d��K4���`���g񔵴�(��	�D@��V4��* ��P��ĭ?m&�$eRي���I^�:쁥T��xc@'<��������[���ۥX���cl/����\�eK����ʬ�����70�k��C8�.����U��%����<yHL:M6�����ޟ;*�(�x$ `���EهPV�ϴ�������?��~��~عx䍦\�_ �Orx����٣��(�t���CX�/�^�P� �[��(��u���5�!�@�4�[��_�����a��42��o�&(Û٪�2�ݯ���a�M:.5�t�=.�E�Gf���X����Iln$�B��77�ƬzSNH�K��b��G�`���`2�+p�-u�-���5X?Ǵ�hb�K.(O���|ntZ��A�|�h ���B�����d~����4��X�_�c&��nZ^�3`Sr`��,5X�
�\� ��eyT������x�3�uᲅ�o,ZT����s/NVʧ�9�Srҋ�333���N㬜�Y����� ���f�\7�+D���X������,;�e�Q��4���q���qrgUڏ1�`�6w��NY3��p#����Ay����g������wʶ�o��e�Mx���8CNe�6��Q,{��ɹ�dkb�d"���^:{�:Q���,vӖ�K;Y�g����FM5\��%���Ү�xI0��y5��4��&t��c��L�Z�^���Vm���#�U�C�
���3CH �����t|7����Gs�p�w��|d���@���/v�tk �Y��.,z�O%�Q�5 ÒYM�4��p��{";5-���@��]qѹݎ����j����#�AGM�Xx��E&�q�!*�	��XD�Pa��]=��G@�tz��E���p9v���E�@�纉�q>F:yAC;�!�Q� a�:Q��N�9�廞V~:��!�4w�Ԑ����h���k����H��v{���X�%��¬�-�̬�GBc���7��g"���и�y`2�p^�E�]��6G�V�۵jCP}�<.����)��M��ݶc$�����\|��p�-Jt��ج���+�b쮷Dd�c���+A��֯ �l<<�Xax��-�U���V�Bk��!��d8[����ET�8J5"��j��5,}
�m�z��aOHx��/�>��s����5���}~^�3�=$���}�v]�"m%�����|�� �R�ug�'��S޲�H�;θ�6�44L���ͻU��"'��ٯ��Vu3���%3u���a�:\��a�,��Fgm³g(4�p������WƼl`����Z�{��>�(��W- 2��y��a�$�XA���q*�^�� �P�r���J��@�Zd}��O!)�˔֏�b�qn�G�&�w���!QQAB�
�;�Q±軲|^�tuu�R�o�9�L����Pd�S��^;?�B�j�g� �X0�R`�F�:3!��c�$�䐙i��������Z��X��<J��_`4�p릛�hG�ͷ"�S#��$�8��Wț�U5:{SJ���7'�Ą�����d�<�<��;%/uS��"?!��=���כ׹ԍh�|fA}�F��
]�5&j�T�h�}9	�1efC��kQ�?܉&U��+#حѝ!t ��C��S����t�),$�cY)"_&�~ä��'B%�Wڽ]�R�W�Y�"���-}Ƭ�v�!TQ	q�� �2�ȉ��p�FgVdvv+M_MM�nZ���|��r:�_�~�nZM49�6E���v��q�]l�-��)�K�p�q�{� Z�&,�w >�{���R]��c�F����VKZ`6�
���0T;j�אڲA�G{�c��ឰl��]�� �������g�����1��G�����uY�HTq�)*Ǉ���:���<ل{0ob���IS���F"�c@C��f/ ��)��p�.$l@BEF ���I%�;�k���c��ǔ�����H_�#w2s;�*��^�Mvn3a�-�x��$�#����9n��hW͂���q�]Y��/`��d�a
L�|�oA��d9������" ��A��!������V����ZƙԞ�.؟�s����>�ӻ-Q�'s1q_&-��**���!���`�O�sp԰ƈ]3��HE�{g(	kvמ����̯��� � M+��`ѓy����y���b�Wn]̻Q��E%�^,���-)�4�N���)���6��o��=J�����NIPo9h��A-�;�W��D)O�����{�4E��Pfzq��}y����7�&'�N
����o�M	\�Ș!��F�h���O�n�VV 6S(��e//w�4����c�&�wR�%떯�?;�A���?;�r�����Mh�<��d�j��f�|���b���ă���gf�����������M;-l@�QQS�555?23�jk���ȈIH�89��ܑ��R�щ��d6w�7;͞b�{�557daQZ�G��W�؞��`��������/���&ɵ�ᢉվ�>�
�L�ё��z��^/nr���(26��^�ǣ�ĕe6{ѿ��2�]{CY��'z�ң�������ҾOвD��wz��f�-_7��Ê;��3V�?�N&�Wm��$�D-�eν�2���v�l�����&� �	��g'�Q���p�t�T�4;�De���.������g�~ee����2~�����Θ��W~��~�/�j���<�������;�a~~��a�H��NL�*+/׷���	����F	DEE�����d���������×bP�&�a<�} \��G8���>6�#5�.��2��}1U	s���g1Il���ث֑�5�^�p`C��2As"~yyQ"�j�����l�����ȋ���3G�N[XUSOO����p0<��9�a_Dg_$*j����T�Gw\.���w�$Q��t��b���)�ѥw�
k��iX�+�z��OE�h%>9���'K3���SX��FM:���*��x��<ɞn�Cg�c����f��1�(��E���|`ҝ��?�$w
iL��b�s�LoK�����`������NAZ��B�g�=z�*�t�|cKS��t�",,���������ol��ﴛ;���@���F�O)�qU�A���k�1.]|�ؓ�+(�a��u����A`2�u��В�m�M6pP1Vvb��=��p��h�r� I����8���69Uo�lj��6x���N��� p�ϒ��.�#4 #��C`�����,q�D�Ǔ��%�|L�K�8'��x�˖��6�t���솛dc3>ٖ�)ݸ��G��J����L�,/�Н�b�=HU������x�cj�c�"�j'|�y�Ʌ�����\�K6�o��G%�7��=����,Lll=�q��2w��ui�--��++ն��33O�W\���:�w�Q���'��F�6��hyQ��zJy1��])(^�>�T������?���������r����C���K�������_3�`��/�.�˝7'K�����p����i�眙�P�R�AP�z'�������,�z���n��[!)��Pjp[3Kj����A���n�IJ=���,6�5��nH�n$m\�ڙ��>���0ӇTV����v��CIO>�VלDi�lt���YZJ���j�~0^��n��&�A��6җ'�d6Ifdb�9�#�e����Y|:�"�eMe�䏬���
	*n�@^�PG�x�&�}�3ְ�@v��~��k]��|��Xl���ɍ��_Uu�'{dtT��������!��kOB◜��M�x޴�3i�w�E�{�#��#�ha�b��(`?�Ob�;�3����k��2�aő\�_����p<I�(��,=y�uT!j1T^���"����/M~cKNK��\�莊��EA��i=j�GǠ����������H���rS3�>e<Ӄn����&���+�jQ^�U�\DP\��K#��ͧ���r�K�H���KVi�J�2ǲ�Žn����v�������+�H3%z@��]@��`C��/]�f{�����ۻ���64�Δ�nj��b��pܡ��J�	��_x1v8x���ZZ�$F]��Ya��ts���=Z�]�	�E%�40���Q���#ml8�6���SU�\�(�p�F
CH��������m�DGG��|<�P�+"�R"�7.J�Wwy��=@�u{l���s�=W�(*+O�������n�U�Ka��^F]�0~bS�*���q{ۊ��ǼQK2_�G�'�XA@�[�iT2����F-�DO;��v�-�;T��~�D�5k1�eN�i#��4i���{��浿q��{"�s��"BC***�O���u��5E��m�r�wx�
x��<����"�Nk�}�:��T��,r���L�$PS05�T��n2��1�Ȝ_�=]d��s`�#EV�nR�o������隝R"��N{�6����B/�ܷ�~:܄�^H(x�f$�
7h�A���o?�^N�b.
����|�4K2�fU$ppp!��RR�SS1� ����{%K𘘝
�����34����������B���YՐ�D� �b�Q�m�>�C��Q��4'$�/++��z�GYϬ@�tK�o�1��eeO�<D�<����d�u�[|�b�w�q����ҿ���f��_Q���(����ʂ�������J�z��m��)oS���tw(%&>	Rtwe�KXe��TŖ����Q�v0��R``�����|�߶�m�u�,ŝɎJ]��R�k��]�����p�Sع��"�ﲡO�.�'-�K����8�2�ke\\_���7���pS�\�;���6�l���# �O�
~����Rwl2�o䵐�����L�¯]F�i=�h�&<��݁�/�F���O>ƋI�R+	@@�8�`��R�r�����%��v�7'}��[�����^��������
[ZZ�=SPP�p��}�TG�-����̆L&�8Z��je?\���ٰ3>�&L>2�7�Ѱ�V�F?<�{>��Ί��q����$$I��g�?�b�e�N�>H���b���&�R��,XUt���~N��o�D	�)��MNN��z����#/읞a��EM-
��F7R�K�T�M�l��syw��q~��>���8��EE)�����'l�� �-V�������p�6VT:���=3=r1~lrv�j
�-�����u�����*��k����h\�j��)R��̗�~4_�2S � 4�T��Y'ԧ??�O=7��@	�n�)�����ǳ�����v��j)������OlD'�?�2�Lo����.�&	x0Q�zF3x/F8ײs�o�P�>�
�%�q+�=��sE�~�M�P* ���"���������?W�}���ol��eק;f���c���f����R&���8�U[W�P��J|A�"�@�9��Чn\��P�������%?�|���;��-��&V�����|D��.4����B�

�.���L+�sw�p����� ܄�f�~����s�#-�[����C#ø��N��of��0�oN�^��~_Ϝ�U��\�V�;fzq��6�bF�����x
"�zW�F��U���	�̰��6>�5wjT���*0�[��	��'����!XH�jo������>������h.����ݻw�pp�>�EDDd�^�Nf�	F��H�Ɔ�Ƞ6Gi�3� (����İ~�!7�,,����-����Z���PV;�H��!5X��hg�ݏi��r��L{2�W����7lã|�w��'GMu�彿;��V�?�kL~6�oI^6�Զ�V�چĒ&mGgg6�ce�)E}��f�i�@��1�Yn�hp`�X�`O�>�ƞ�7�"5%�x�X�:p��b�C(�H�H2jo���e���fy���gV-ԫм���������@�憁�K�nV�ӏ�<��'B������i8��	�R�i85U�?3q9c_�}	�T~2�2���G��+�{�
���\8��g0U [Nh�������j��끭qy63W�T�_=��k5�o|�P$��==t�tm-�޸ �r��Q�	����Eu>}��RTPGFnh_�RUQY_���r='�q9��|�8�.\�����n���A��ި������Y��Oo
䳢�v��i`⬏S���Ҷ�`N����3�lV�BNei�
Bű�O�:G�����08��ۅ�"��v*2����Fvt�4V�T�ՠ�E�ܓ�7����ON6�cy�#5���� ���8�=%�k$� e6�����nk:���+ˊ�*��#K��5��E�J34�k��R����)��:���z��0� f3&��M�#�������i���w���s�ooi�֒�-�����T�3��|)-�m��YcK\[�.�#5����%^ws�1x"ʊ���Â��v.7F 1�}�R@Kf&����LG����r�? 5�����z1aڷ=�e����4@д��*|̭mť6ss�`���QT'�*q���m��D�|}���ۊ,������@6�Y�������Ն��i߈���HQg[G�>��� �"�K��qUm����h����Q^��d���]���.�7o��ǁ�~�7,�|e���;{J�4?|U��Р��g��D>�T_�A���	s⎪־9����79�$Gx�������Ĳ[r������\��.BE�8��<VA�qqteC�Y�El8Fi�3;�����x=���ό�I�׶7�B���Hy�P�0?VVa	���PX�����L$�P<�3$\�=S$4�WT�{�!����ٜ�]����g��	�ɺ�����$���W�{uK��G���}�i��?��O[�`�_B�����F���:ٶ���w�٪�ɲ^8?���ۛ�>� �onN,���z>�44�]��:ADr���I�lk_�Q�*����t��ʏ��H[)�N�!��k/{�����/|��%��������3�߽���.�d�*�'A���!��iL����x(��)#�w�<P�ﱰ���Eȓ5Ry�S:�Jy�E�G~����0���Pe �%�e��$��\�n[��C��a��)8�QEJ���}5�Y�`^��n�����^�v�>(.��8Zm�(kn1Ԟ%��S�U6�4/79�y����%G$XJ����Ε��n��k�h��z�x]������T�Y����	{
2����RI	؁���a�݋7@����
>�^3���k`@��Mb\���\����Ͽ;�rBx
 V*S���17��ۀaC����?�j�Y�2�n 8����*ժ�
�F�2����X�f��ΐ�8㕴�'%Q/ބ�WB&�h��Բ���5�\��8`g���O���a&&&\oW\�>|(>�&VY&��$��&&&1[m����^�M�=8<�T`���}E�/�D�߰|��{�<��5x*�8�3�<[��߳|��f�
F�����a����g��l
�|�5�FEG����c_b���v��Ѹ��QGMYvN����HM�������R�y�]�������r$��� ����Y/�GFLZ�V��r���¯�,���"*Q1����do�֚����iU\���a]Y�000���q�F%juC%�V�1'4��~��� h� %ж�3��#��]`����!:!mm�y�w#��[7%���ʇ/=&Q��1H�����p�[]S���E���ӭ�N+��>Y�O_���	��_�5�尋����f�?N��wB���ܪF^>:2��!G7�![iI;!+%e��vS�8Py����b켷@V�H')�D4a�_�z��-9�2�BAr��=U��U�I��L���cH;\��妓���8�̖��Iu��9���;W���V?�����G��O-"��u�<֢�tC.KJx�Z���E��I�+�ޢ5d~�������j�������E�����Hqb,���Ş���B�Ԃ�^�u����Wx��c{8����
�t���+�e�"���G=K2�p.������KK��i�v�z����,o@ >���a2S3Qmy��,E�C2���s�`����Ȁq�pllm��{�31)��"�2(2	�p�~Ep~?$���'�BE��i5^��ۏOj�Z�j�sý��iq�~�S�	7�?�(�X�(1��F��F�j�6U��H���+�l��lmm��`͞f�)����b��x�b�0�3�����K3@��Ĕ��B�)�c���Iay'�H�&��m��\�u�(���G����t�8�S�H�zMҸ���W��"���D�S@�4�^|���ʫ	�}w��F!���E��G�g�[����}6\q��O(��p���U���B�2x����z�4A���0�*�'T)w\ߚM:��y��5	�~���]@M���v���|#k���7�����R:�<�!��і*
�������Wt���w���	��=g�����L����{xXf���b D�����fP^\ѻ����\ЏS(_��X���' �T���/����*��'�H�j�F����H�0��hzf̽7b�kkD)))���J�\�wLA(Da
p~���4����C��|n5��x��=�b�Ę���7�ݔD�^����v��;g��BON�/O��gѵl�d�2�666r����U]`����B
|		�)lf� }P8�v�À13����8��b)f�x��������t��x����w�!���q[����ܖ�{8����Z���U̍qb��
s���=T�GR�)������Mp�Vʂ���놅���NK+9������]X�Z4������g�mJ�Y�X�2�Lf�,������#�Q�Q4��<7�1Q��Fp4�� ��;^�Q8mVrr�㶴���=n�Q)���QZR+O���W���"�!r��9�tW���0y�������FL�`�`�"���|��� ���:6���������dB.(���z()Yz	%��J�C#%��b~8a!�ҁU�F��b�h�F��
t�o}����'���L!��X���iT�I뮯k��,W���>��\���b��@铴t逝r�\��P�@zp���D�A$,>}�ۀ�$9����3�3�|���`���]���#�w�����T+FL8���EG��^w<������}����j#B^ъ<��3����������4-�����
*�:�<�p9��ҽ����:6�c}��15�V��d�=:�U���ƑK�?2��x��*l����/�ߣ`�܈���6}��ES��&��������
��˵nB�h���^�?��0N�Gvm����n�r�ZT,�v���پq�-3Qu{7)#����ى�h���|-F>b���'��n����se:���aU�R�Ɨ����>��z*�r�k@����E�]�s�KH�HD��FGG����+�-%��k���f�F�Q�����`������E*T�}�XJG\�{�C�&SiPr����v"cV�n��ͩ�����B��$����l���K�ӳ�x�_k��ܯ�\��]΢������3X)�ѯ�����,�h�X)Bf��n�M��7NO�VZ\��0ppBȥ��sD`�������R����\7tJ���� cnnm]UvԷ|��"�셼.�ϼ2,��7�ж�FP�b+1�:b�0cJR�j:0�V�z9��U��8�)*����#�A���C���.��H���3���0^��H/��"�Sp��p옲�M$��P�N�o�r��,�UuO�`&����w�I�T �g+�F7'�}�W����0��?,.AES.�dN=H��4n�9�	�[�x�Nˮ���\Z����������p^h,�ԛ$�[QQI��M�O�SR�⿭$�bC�z�6��^��;7;;[���%�|i�A��^'Ve�L.�������;�\��bB~w(~�6�~P1����������/�I��D�Z��A�_?���t��T��{������U+�<�*��ॉRox�'CK�ptZ/�[����_Y�����l��w<_I���R�F^60��_~�1��Wn��������+(��a�Z�#~����j�F���,���@!���C�������)�	j5-��'��x�������3mk8U�Ü��y���I);4,y3�zQ��9{L�R�����ܸ�HL1t�_��Fr�m���M����Lo�6�f""y:��&A�Z��݈V����Q���=<��5d-���b����N��5_>f�k觧������جP�'��pQİu�R]+33�|^�z����eӿ�13���y�kk��ze���ܝ��_�N�9^膬��6�]+̷|������Υ'*$����h�4��X�x��t=�+�xtp�4[�q��?{����Q�Ȉ��]���^�޾��F����Z�%���V�Օ�B.=�E,���n��ǿ�|����lǆ�����Th��]\\��)��%tJ [��P)����h���<_�D��*�7ʋtτ���	���8�ґa�����+n"�FJd�՟�ҹ7>3�1�]8�6xHBM�y3�DG-����p֤�l)�'���>�����`���Nf�!1ssB�m��Tiu�5�n�"^�&��������٥�~Y�e�H�F��j��I�W�'r���;υ��M��%��e��:��=�(�0<]�ZD*����g\��H�27F�-�j�ʆ�]���tޫYE��[Fn��@b`h��	cb���Q8�{x0s�9/Ez�F�S�^�i�3��?�������~ �$L��3ɌV*�)~�>���n�=ug�����ײ�Y�][�RT^*�.Μ)0�WcS��u��|A��,� OM��n����L�"�X*jjaVi���t���P�~���e��h���o����*�`�߭��N��L�a�T�����-��r�b�S��k[��:;;��@͹��>36���juUT$�:`�1]���y���0*��AҼ� bw8�?����L��z�#5��������8�'sXiִ��!���㕡�������1���ur�=����m�Rէ�q�䀷��ݥ�}���&&�RaE�[mn�F��['|�լq����^'��U�Fo�71)����t��-�)��/�i`@�5�E�aS"��8u6�G�m��ՠr���Z�9��U���[ZE0y�0�*�O���{���<�>F ��Ϭ(�NԏD�G����-[�w�g�1�<Z�Z��:��Cח�}>S ����[Ugɓ�Ԇ+v���䚪��m}~�EǱ��F���K�"�U��_������%��o��%��f�&r_ԡo��eύ�3�H��\��-w.a��s�~/qd�o\��(vMk�N=��i��Z�,��c#_o�[:���#�����1����F��Q�LJ�C�n�|}�"08�i�E(���wJ0��u)�\CKm��oC���5�[i��R��;G���Ӎܪ�/j3���I�^�}r�N%d0�M��T���̾�DVX׷�����}�JZ�=�8=�����b�7$<2n��~�����1bT�	pq��w�RB�=?\��8[�J9`bamN���yܢ����X�n!�騊��n=�*�)
!wwh��؏1�،: ���v�G��X��jC%%�x��.�-a}���tt_��X���A�+r.y��9�B�˞���s�u5a=�}�	�E=O�IW�:"���^��3$W�����ߏ��n�t{!���j/F���
�ͺ�|�n':F�hI��7�����o��֯�%��f{�����:ս׮�9%FϠ,�������ҝ�<&�+�ږ	#YA���Y#���_^��
��U�8���k$.U�g^����搪�6�C��^�ί2Q�O�`|���\/�2W�i��V�a,鼫�u���Q��a�M�َzKTH�t�`�_���&����m`uLT�%F�uW��"�3	���G�[�U�D�Û������.���i)I	)AZ��A:�S:�A�w�s�����|`�'f�o̬Y���5�w���5V����O54����<�%�ݓ(��bR�v{�<����g,����QKvvv?
y�����b�s�ܬ,�S
�	����c��,,�������q;�R��{�����<�7	���ܺ]�R�X`�3���a��ɕ�Q�`ɻ9��������ZK8��(�ꀿ��52Y��h"h�\��������P>��~vvD�m9 ��QS��^��u�;���k�B��&ИZ���Loޡ8��c�	����a�����C4y���񗳋����jq��
͐�2)ё�V�/K�������C?����-�k��a�g�~����*�y��A����h�gy�v�G��9��,?�����W��4��)l�S����!��Ah�o��L�J��&��FQ(qjx�0��t�����cmn��G�/���-�1C������o_��T�R}r,�������x����/Z|��&��!=m	jr��RC�D��i�{�_R{aR���9�hĔ�O�juu]s��%UV�`bRN2�ImN�j(�}M�FK3!+�B���&�_-J�H�P�J��R���[(iN�¡���_�����}�h�mVs$�UC��vQM �

I��F3xs�o<��9)��:�9bWǿؼ� � ��ml�TrDѣ�(o����d�((*ڜ.Q�#����I\�D��n&��l���T��F����G����^X���K\�.��J� \�|��vf*9BUghs	�q����~������&�jx 8�uF[��TC��ߺ��h�ŝ����������6<X)���Wx���ߏ�LʦK�^��r^!*�gA�h@�,i�[qZ;{�J�[
~��L�e����{	8a=�o;��UU��!����4�>���lh�pO1�r��M��0�jǈ*!��s7�m$������a�!���x�4>�.�d�6���Cv���<ݜ�UgN��H�_"/sf����$�`�+��f�I�X���̬������M�:>>&�w|���J��;;;Ɯd��"�o������
����pJm����̴���wt��\C)�D)�Mޯ�xG0��'��M<K�yS�5ݚJ>���#�[�Pg���=C�7�w�N�&=Bo,oF���K��s�����1��T�ZC��Uo�v�bﴬo�	NO�fޖ`!�SrEG�O1b�Y��n��m���ؾ�"�}�^��mdTyn�P1���H�Ȉ��/�J��͙ށ�k�YʯÇ��pR�
��ۖ-���j�-�z_��ԗ�d�?������k{�n%�L.�+��zY�s
��\��mM��ۈn�Q��E�=[���g����@7�2���(���2��ٿ�b�W�W���G��ЄCƃ��,���eS���(D\f��]�$z�s����/��>��Χ����k�"��?'L�K�rcS���ڜy�
]�<�?��E�B�@�N��	������wu~� WR\��BXW��1�3��W���uqz�lS󟞆��Ɵ0��,������Ǹ�t����T�'�k+������qjV�z�x73�KaFF�Y��,��qb�ק���ιzs�%~#��J� ���,�L�����3�YcF�Q��o+��9�gL�r6_I������%����w��Ԍ��;V��^$�|U{�;U�D�>��^r$����F��fƎc�ދ�v��f������w�8۹�ȸq�+��K���z�}����e|�<����-ډ�]��V*p����U��x��{I����X�`�퀊�b �ҕ�Q���8����7ӓ_�ي
�b������U�~��8ZXX�>͝o0	i3���an�,(��S�q?a�����V�c�G9_I2�/�0�;>9�*!z���}HHf��D>
dЁxj�NF�MH7�iC�x�M1R-<w�eMI��Ku2]�4}n���ֽ�p�	%hrRf}1�G�򵅅E��P�L���8%&&����
���\{�j��PA==vp�$��[}���*$k�G*�f7Z����Ʉm!8��W^���0�
[�0�~��樐?��-��o�*M��T8��Y�-:3������A�6FHx}�2&F��7�qz�]$�x��P�3?���B�� �/L��t����n%x�o~iy���|��1+fH�|�2B�r�Q��5&�X���9|iN����I�8��V�3���	
�SC�Qb�7]\���>�{��Q˞_�(���Q��%(C+���֏�7Y�PXn���tn~����(�u�x!�v!_���{x�����W(�ty��W�������S��� �D��� MR�y��~�\W0�	C�;�&��K�D���E5�[��=������M.��o��OV([Z�襓�x]�H`�SE*p<��j%��w��F=�wz�C��g�)Y�?_������OYk�4'Yx�0���5���K�p��v�L&�0��F�:w�m�aRcR���p�A�i �c��;JI.���^����%۹�x�"6�<��TLb��ޅ�&��j5S� �I����%�~$鍇t5+�P��}�D2�	����&n6�:�F悑W����o�Q ��ǈBє���e�QO�������5����LX����~�ެ�c&zO��B{�d5���L�RN��h��atu���F��W�2��7=��FN ��?U�k��9�&f�t�|�����øZ'O����P(���������޿�*P;�xXPFYo_�����a�`P�0)~,Ñ����!�9�=6�!�+�����y��7�Q�P}���ccF���Şg�7I��Ԫ��{|�3�9��tM��T�y{&�˿KD�|H��LIQ�I̍��З�~�:A���b-58$��_ [�e��ò�Ĭ�Ak��T^^�x��u��tSgzzz��b����.[x�r�w���FW:喡u����K�����t�0)��$�pa��膅[���KEﮍ�8��"z�׀�_K��VD������ns��G41�� 	��Ϩd���J�ςn�@����B]��)+&��գS�����_�m�_�~�	u�������?�Y��,R���	��7�pqr2Q覩�*���lq:
Yȗ����s��
qsD��~�D�wz*ay�eO���:U�r�FFFM�ͼ���1%�qs��_WG���k׹zF�(�9��0�=g/���tn��Z��w\~%!�!��)&=#�{l[2�k ����x��;��L:�X��ɓ���Of�q�U55�%�EP%��+m~P���?��E�L�LPQQa���;�����*�jK��c��.&;[q��Ƿ
���l�P�S\�$#K_(T�!x]���.x�Z������h�)չ���s ��Tӄ<Xg��3��0���U:y�8�' $���#jt����6����P)3|"_&�n���6T��������'44������ǻ����� OOO�h1A�E^A���Ԙ�'f2|�h_����bQ���`��B���"/�T)Ԧ"��˩��/�����ǧ��|������5g����]��bf���D;'�}M[{{�\s�6�2�����R�9�ƒ'XV��+(I�Z:z$�ϝ�����2B!L��dC{"p̎���E߮�y���$�+W
x�������7p��8�=����(�-�� ���Z��rݐ�������JLNxt��)��j�>eg�z�
o�"vO �f�!>:�'�^��mW9�o�R�ӪhhDd����2�.h�V\��U�S�ǁ�rG�Q؛�+{p�p�o�(=�WX�]ɧ��LF�u45\��HB^��OR�Tk���v>VLȫ�zbevD6{�D��i�VJq���G�(�� �$UTp455�Q�{±zfʴ��\&�sM�>=�||0]��o��O/_�,���"���Xnv[__Γ���c����e�j�ښ1"
J��L�K����� ���6-??1�$	i��͖�:h[�N�7����D�����n�e~U.@Y�CR �� m}��kd<j��s�Fķ���X1Xۢ*��u������_�FW�Ȼ�pr�ż�,�������f�$$�ư���-�R���j�rE�'|||���*י����!Q��Gg�����U��_�8�8� �J��7��p�,~P'rv���_{�]�/����L��Fp[�����������++�NL�GE���;opqu}�����*OUUS3,9� pG�0ç�j.a++������Htuu#��#d��?�aY���;99�/,���Y�����P��,�TS�O��S����:���@͋��V�)S�Ѽ�������-SQ=�:�p�:�F�}L���������-"����u��АN�ޱ'���)��Җ
}))�B����#��ɩ�N�77�_��>{� ��B��i/*��@.	:���E]}�� s���S�C��f<����ju��82	�������_�-͞qp8�=a#�����S	~�K����a.�C��_ �3��_߉�����j������������&&))y���JF�6�����ۏ'�p����BP`���?���'��6�\�����LME���ע�23���B�={@��񃪽��Vb �i�`��ܤ�;Q*g�SSS�0����;�w#�/� �g��U�B	������9b^�8�,��a���S{��S�R{��Tv�IS#@v�߾������t��v� �_�c�)sT����L�������!�1��V*�GضvvP���^)�8������C�n;�N�����t	� ẁ�q9ߒk����2J����B����=������)-�k9P�h�ᾣ�B�T�TNX&�DGr� z������'�ť9�!�ަcaA�0�q#ʊP�g�������{����~T���d^:;F����߼@���#*���(6 `U�ef���E��Fvus�A�"��9��^���`eeU�����Պi7�tE��Q~Y9�.����.`��d��񙚚B��D���*K�X����T��0џ�3e �N�#��DE��rNM�*� K�ғ�ξyoo�sd�{ 5<"�p� ��~�
>��=�����М���(���p��P�S�-Ԛ�hc�-�-�a�w��^=ssڿoC$���l >7j_�Va�ߥ�����@�[c1|��k��A����dd���	ֻ[T��?i�����&��`|�Qʞ; }K��T$$��[5Gs��ǉGr�l\)W� �7M"��D�����������1�A�zx`�@�w� �IThA��!PVٰ����:`�X��T��)���`�Wf��LA��a���,��U|���7�Z��,!�����[(YaX�
��QSs��W2_C�!�v���g��.7l��~������s���j{,P�t��E��*<���P��Z�1g��/���%��VV�	 UBG�����p=7h	��2' &�2���CA�q��WΟ�J2��"�mw9����
*�ꏧ��c�ߔ��3��-[��M�ϧ�v�3�A���=�����7�]�Ue��ˏ��:1l�y��2�����" p���I�;⎻s�;�AS���h{���`qEEx^mkk+���H�t\R�(����Wv�D��"ﱬ���[v�1�'�K8��춛�����(0���X}���.�؄�*]������x� �v�ZZ�xv�a����0�F�E�B.!I��R7}�IHw�ףsT�*&����O�X�Dr�@��� �O<�t�Vg�9V���������O��{�����+(@a`�Wekii���Ƶ�0g��/��Z2�~�����2
��2$H�h�ǜV����_-!��8A�[k v�|}��Y �X�>}���.D���H��F���oK���_x1�70k�&��OF���]hv+ҩ��Z��K�� -/���14��3�C�gO����m�z��wg4����v	I��*�k�G��;�]���k ��\t���S�N��R\������
�]�d''�Ǉ�	 �О�'��������[�à ��^e>��7q�m9�
�y/�J��]�����ԕ�1���l�wwg2솭$����p�hih^��,��Ti��ņ��6Cc~M�{��Q�9�9�z�$v(1���ſ=����R+�"̣�z��ɷ����?�]U�kz�4,�:�6a̹X���V�2�?hԑ:�Xm�B�qy�3��M�_�<�|+?\g�@'�ǲ����u���v��]-��ʓ�$�1�bT�N0z�ੜ��J�����`�������Xa�0)�;l�n>�3�m��.���9<��q�o������Z��z1���Ŷ��Sʳ�[���˨�7B��wx�O�л�z��7--,D�H��X,P��g�`�]H����p!(������G ��'+"a}��D�A		x0��ϱ�M����a�[I*� ���z:;a@�����<s>]�v�Â����	2'�d�@^���84�U������g��돵Âu�wszԸ��hjJ�I��վ�ۛ��?{o���X�������O���k�V�(��KT�!>5��e��2ς���`�o�C�L}����eV�O�-+z��A)��O�W�Z3_	���|���c�Ҝ�h������_UC��kb��va���\�OM�y~��׍ �~t��.r �j����V�'������Q�;�QV�%�p����#FGF���C�9�Gx}���� 	�w�WG�_�|���^&n<5�cf���� ���=�$U��5 �{".��YYY��m%��ħ�i�Ð�)"��7�m6~�i�������ٳguN��#܉T>>>���Vk٤"/$�a#�+I+��"47Dj�jh�3S�@$9���e��-�ң�����A9q��j2["����I}�!D�F%���T�ʊ�T�$<s�s�Tja� 6튵�L���m -sKJ�DDD�_�ZX E@Ƅ��6����˫D�<Z�)�v����V�E
�Q�� Ӵ�_�ɚxzxx����'�hށK^?��`	{Q�*��bM��$�"g�6ɡOZg��3KP���B�|�Z�|�F������^P�@L'nC�!�kq���K|��-x��m�s��U����L���"��;?�VV@�l�C�e���EDXp�{�T���S�aO,L�ys
@�?�ƀ�Eƺפ�˗�?���-�U��L��g~���G�ɕ��eǤ5�b�h։�֭���\����"�t�\F!+�]3B�<�h:��N����7��i��O�>ge-�͞ۆ���F��x�b���yՓ㿫��Ȉ�������J4I������g�f�V��b��H\s�Ͽ��nd��ݥ $d����or�'��@�$	Zjt���d("�T��݋�����t$�� 	YY�@<�rp�XXXx�^=�:Y�w�����*G�u��^7	z�@���r{ 9��+ ��VD75	$''Ӏ/@BB�~�y��{��TQ�A&�� l��Á� & �����/�|.,�nU8ԢR�����
�""��ZgpUCӠ%p�O�2k�i��"8����i�����5!���abp�'��t"�l���j��NO��8�hZ���r|��9�k�wu�x���@?�����49v�?a]U_�C��'���d����kp55��w*�� mq���9��Sߞ�6�tp��Ow���2���lìGff�M`���g��p����Π��ˮ�U��O!�&�@��tv落�!/-�9T��҄���	j�0:��K�?�2�c��"��/5�y�k'���l�@�WG��>�  ����{m�����<��i\f�߾=���+���r֑�w�O��j�!V�G��rsYVkO%2o.ww6�SYRb��6--�9%?	YOO�8	�#��7�Fc������._"��X2��nLᦖ���"��5�mw
JJ<\�γ���RVҞ��\�����[��spp iX{��Ԑ�kG� �m�X�q������
�y��������s���A^���iU���������o�M��Q�n�1;�M����??w�$�|e����D��Q���Ae�<O���L -�-������ޱn��*�4� ����"%��������J�7�p zY_2��Yv�#���m��~������s�����B�>ȴ��CT������q))G�&���������$�4㖶�n\�i��x;;�7��<�m~�оS��h�v[F��`MC�U��P���pQf�ms�l��㲲2h��q@@��J���%���f�/���������)~(\Aaz�?#�����?�검&�������CX3������6WE !���x5�^ ���?�6��xk����m:��@���`������ؘǬ�H:���i�_7��׷�=x ��r�6�ff��.�|����P����0��u [{ ֓p��Ar�&�W76�� �K|�u�v���jUc҃���"�ߵ�jD7����߰��捪�����@��13��qy���Q4p ��@K{{��GT����y;	�"B*�����Up#ͥb���ő�d��	~?��9y��׎�9��rOP�ݕj_1D�d$ͭȯ���:24d�s���8���"��Xl�e�I��֔��!?�gG�6%���O�̖Hx�q��?���5p������B�{A>;�BBd\\\Rb�M��#��L�В�a�ˢը��㴟�l_�����a���c�����t�{<)7r�t,��ȴ0�g�;�Q�� g��EACCß	����H�i��W3�����J�8
A:g&{��\pA�2=��2[��!�E�ET	d*�����!����P�K����G��#��Ճ�.BZZ6��	�-fff �����`'���$
��K�||ȝ�|s���s�teYĔ/={�O�c�6��0�!�|��/��*��s"[%����@h�GN.f�V��r��+�������..�(2�
X��} ���u��ݑ�����e�TB������͌� ?p��<�&|}���x������pk�W�p
/ٷ�F�;A��?�폘�H������`z�ݗ��@�J|�Ѡ��u$;�{�s	�ׯ_[��~h��U�щ�<x}?�������Y��A9���$-!/S$��vv�.9��R�s�O�<�AW::�H�>��]���Zl��7�onJ�X���Gr,\P�_�	�&��p+��Zr�34�n_ܧo�H�#�ǆ6p��]�����j�Cy�1�L��H��9x_iJW�bb9��]f�uM�88 X�.���O�oѓ��cG}��9E����˲xOO��9��u��x���@�+D����Ξ�JO��-�졣���o�_x��;�:�����n�"�to����9/77�������	˵�V;�N���\��cjrRjQ䋜�	�%����S���f�N��S�i%T�ӗ)�ʕ�a��49є	ޱ=~�Q���-(6��8H����q}�M�8[�7��sv�ү�i����o?xq�ӡ��L�33x��j�w��U�������j}ӃN��漀X��`���{��<���4��:dY%%h�O��c14A���ka������[��	�N�G�i�/F7R��`��\<�--E����`D*�Q��Mנ�S���8iii��!���V�ǔ
�T�9�x������! ����/t<<<5QQhK�k�3T��hlle�C��,��8b_>��@|ch�͚�rq�{i��I��OO�+4������j���'�����<�S@tV��_����כ�b����\�c�p����61o�B����c�����a��t2�\"�7}E�&y�H�ٹ�@W~f}��o_��_"���	�ou���:�ǿ� `a�l���9�ņ�n`|�ʯ-��hbb�Q�C��u|�&�2dc0*&fo�\�O ����P		c��&�7~��sn�������l�:�d���k�?��$;�x���~8���� #��^��:j�8���mm��V�<�vvv�g�>�>��~�j���z���`����L-�ͪ�XalVi����J��l�5	�yB9*pz�F7�۝�6�g7-Drઐ�2�AzI�eI���2���g�+$!�Օ<�	���t\쑇\0�������F��
'��3<��q�X���M�!�	 �Y7������0�q���䔔�dEa`f�>����a�����"%�_MU�]k"�]�J#�<3�7^NZr���V�&
+X=T�)E�[Z6�������YiKx�l#fhD�v,�lBEq.���a�,���w�G��h�����}}�==&&&��ֿZx�YR�|t |vu�k).+��P��1��%mpZ�S�M�����s�J��R4�O
�=0�q����ӝ��@�/!��-����Y� P������+��ꕃX@:ou$h\�>��B�A�.������b�0�>�pީ$����`�R��߿��=G�rm_����d%(]�"5���`	�U�KO��<�6ߔM���Bd �u��a�n-@�!Rw������㯦�t'~��N���w�T54
�')�`���ק&��=}��!�y�x))��� L�����"�L~��
�֐�CN��:��5 �㚸�nnЉ��vFFdj��g=ݵ��x�����;t��޾��!?222Pe�0�N��������>l��~����nle�/������?��߄ �zf���7��&�����}~~��L��Ќ�������UUUA�C��	��Q{{�¾"w����!����T"�?�u�p�����#[˸�֚-?����{� ۀ��ˣu��x����L ��^PP�:�jy��ʎ����o�;��F�T߼71��.[������Z3v����8��S����V(���'���Ņ�
��O�5�^�<|�0"{�A���c���!� ���[[�M8���g���h���t�,S>6#l.rVCY�-�C�U�K�PYl��nZ�2!ɿ�55�}��pim-�~#.^��������cNcATL��>(z<_M�M-:R�����`nYY4gy��c9b�����><�qk���C\S3E�@�q|��f|2�'L�4���"���z/��Ь,JE%���"��4�`v~iAR�R`2|��{��%A����B1D8�
��G	5Mڍ������8r����2j-�1$@T�z}�]\\�kC
�/��[�O���pf��$7�3�z��R=s�?�p�*��*����3�G9ĊJ�L�dc�e׃2�L�n�����x���l0m��ǭ�����toN�� �wdLL�t�z��Z�L�BEq���z�L����2N�����s0¿ĝ��a����\6�66ޗ��ȵ�}��u����u�靈�,����+k��I�,=��e�Y
��L@d����{�\.�2���y��
9-���@����=�5?��F6���ɓ'ЦB�7o��?��6q.��Q<�u��ٛ@ �h�אk�g���2�v��{/��T��&$�{�TU�����a��n��vF�3�F}�X䲼4�P�?���J��h^5�� �xv��&����s��No���|M]�]@���S�Х�P
.��0J-�d�c܀N�)���XAq1*����/�Z����300�
�z��Ѱ����<!N�F��7��J4X%$$ ]���(B�ؕ�p>�_-���²���9�^)\�̔kw3J��������O�{ވ�G�񶅻��c����V�P3�h�ba�?yrXD�nej�	p��M�����8_����y�B�>	���E�Ç�1N��& b��z"p"""P�@ʦ,K�����/�4Vʔ������3n�-Yo??�l���JJ�<��U򲼡�b�
���ިw�����W.l�XX����Z4��������s�����>$Ƃ�7����<��"�abXr���jH"��A���<�x��:�Z���-��M �n--���
��(Y��ȿ{�n˷�a�/��N�K�QZ�W��
�,�n����mrx-���C�6���V)�?S�x���s>��&�4~�L|dmP@�t����,�����j��d��ˋ���PUU}ec�Z���w�#0�N9#3����^�ܝ�˥����c���II�Y�Ȏ��X�_ժn=A��,a``�QQ�B���a���u������'{��#y&**�����~���c����bagfz���p�M��s^y9f{{;B�D�5
��֨��Ҁ���o��a�/(IHK��ov�e�'m�Afzz�����|��9�����(j:�1EΛ�
=8������~¬ͨ&t�ᖐ�<0'j�>�c��x���&��y����\��������\\
���'��?~ ��˶��~;'����E���f��P1�'���p�Z2����br����C\�Z�Yb���p�{�-jD��jL��������h��������l���SV@������C�Ğ�n2�v�<[m��uMR���P�T��CA˕�<=�~��<LI����#)ГL�YJ>!#���ɪ�ȸ���^���~�����ݽ����}w����� A�����߹��J�������<����3�� i�6uUU�����vR22�����G6��V�����'{{{#[����3�ă�n\�&&f���H:7�7���z���e�"�y(������/��#m��`�)((CƋnP�c��HZ�ݷ�]A�� �%���W;�?�A55|6���\f}�;�PO�R�2��("�{�j���݅���R���DS���������i�,#'�bW'�*d���T�������HILJ��v�EE?��%�Ń�ٵ>�ļ)+)隙I�u#�,N�pw��,�E�%� �����.�G	U��P�e/��x��a`b� ��G������x `n��QQi]�vFֽ)?2��[��]�6
��@N5���=6��X�7@�` �3����1��PWt���Uŧl�P��鲚 MlEy{���:fZde�*�if��J��q�>R#�������qh�)�J���~@?��2gyV���ɘ�iTRQ�sëUi������BmQ\����r�T�3���4�+���1���R22�g,db@�2`{���mtZ�1����"���N`�`���r� AQ�	��*f	���H�YB�d�������[HH�Ös�Z	���d(�Vn�����pA�B�BB��fo�*KK7��	#����vj��F�,6� Mr�J���;��O(0 ��4�9�D�mi��e
�����f������������0�rhz`�qS�c{�g�r�W0I��`D	}�@&��`{�h�|��V����O�Ku�� �ww-^'�5��g�.����y�X㡵9 sN//�jk��Ӽ�F�:��ϭ�w�*���˥(3���]pWZ<0���)�)kkk�ww#>��t��l�������!!B^ǘAUiI�%--dV�ٯ--����h88�A$o��Z��Ƞ0+_ؕ�}O5n4����� �Tꤧ���=7jgO��2�!!#���1絠�Dف��A�D�Z������lI%��	��0�@f
.~<(�:f���(z3`5P10��:RRR�n����@[���
�-�rXf����$ �J���ϟВ����˿?#@EQ��: 2P�Ѯ����t���:�a�EnG��7�::�@�2)e���H�W䆄��F�;"�_�~e�sc�%��g(�LK��t+v�P��hJ_�MhyxHʫi�Z�7����Іn�x��ʾ�EhNZ�������7W44A�6��<���z��[^Qwy0�	l?C��w/�Ո��������["v��̶���k��f>��t�w�+�M�?�0�X2Ə��@:��܃� ����=�x�;=u�*��}�2s4odq^=����su5�=�Bp0V��˗/��M�\M'�r22Н����3�ԋ�S"[S��Em�0�Eg�ɍ��|�dd�����C��?𙐾��<���B�$�4te�5�p"���2A*�߉*}s���?��*-�_�2X����u��i�I��ǌ���؛��7������C�S�BT�ZZI�*!O�9jB��7�ζ��KN	�Ӏ���t唔~�>Ӈq�0�d����f���@[���h���Y���K�;���80<�D�NZYXĚg������C~��$I��/��l�Z�K:��Y�0��)��}VAt
=M�C5�%� 5�FFG��lB�X�H��w��ɈAl_��>�� -6z����������ن��d�m���Ų��T;��=ɹ4a}p�Cj��0	?�f��,��<6L�Җ��L4�u�G3��!���:߶�'�_��0�Q�6faii��f.Bn�����.H��K!'	�s�ַ�
���D���h�	�6�9=��aO���[�|���V����46�WS�{�'&�X�\�'��\/A``a�l�rqa��_+�`�kq�����n>�/2��47#h�e`@���`�t�T+x�"� ��7%4}P��� �.1�`V�P��Å�#��j�mp�[z���L��,�> �I;��إ�n��%��yC�fڍtn�^�h�!^�߼����±o�~��wo().�U��?�QQ���	c�,�C&� ��,lS��
���͍�H����9K��N{ n��9L.x���JR�u��z��z���G�Rے��^�����@~A�hjB������)��Q�֡�?1��+��[롺&��T��������L'�HSS3��~������frJ
�.����m7P"O�ͦ��l�-68dv�8EEEAmm`�u�,pehƲ^F��(.-=��=8*U9??�ܽ�B)�r�%�爙��.ɝ����j�$	"2���>9###PDM�7���\����X�x��
J00�?6m���������J���@���&f*��++��UUC�CpkZ�Z���Ū	8r�H���oo,�m���?|������s`_L���7���U�%T�@/S3�)�o2�V����ID��}4�����
�'4<|�(����������������V+ˇ��v�QQh�߾A��0cs�9~I=ίi����?��?�Wc���l��T�l�%#��^�����ۏ>�込F�<UDG#���RUCCCo�1De@��:���Tt��*>�Ep�%T�oxx]W�Pa薏s��d��p##�+�8���˖iW��kx<"������O�Ww�#-U����h���1�@/̍���
F�&'��8.��F�Oޜ�g�P11;�+J�%tɻ�p�;�p�Y��dA���d����4�Jv�А��[ŕ�g��߇�������~^_�׮�����.���`h�q��Sd,9������~����j�s��O�"Lz�M~�x�6/{4hkht���Sq`��8p�����%H�<�e@'\`��j׬X�eI�Q<�ֱIJJ�̎�^���Gquu�܍���+u�ͷ��pӓ�6	���hf�Q�}���{b99��,{zs`J
N�?�� LC�W�	����x����`�r~���8AV�١�jp�'�����~�{qtJX3}̩�d4��M�s��(��p�3fʴk�e�ӸBx�M����fn>��Ή�^�,eEE���ֵ��X|���)�޾��m�N/�v ���[q�C�����/�����S���3'9�~�<2�n�� 1�\�6��{K�)�����uvsq<{�$�#�H��tb��89_ihd�	����8_�(U(��;�6�M$:��޷���:�]���g�~������-pȧT�Њ%Ժ��)�n	^��(YCg?_ck�/1  �	�/r�zZCqL@�? �W�қ|��or���x��?г���4�����������C�,��	� no�aN,M�(�k���3:������;>>~$��ݱ,�L7��;3 ���~�w4�V �O�q$++�	4H����kGU��I�x�ZV/������#�3*�� %�6��?���2B��Z�����5�Z��5evvV"���H����˰�v�l�x2Z��Z�j&]3s�F*}������er��H@Tɀ�! $�#%��
�i-T*H�[p�&����f`��~�t�
H4�7/�������tDf����0���d۟+�3M&���j���6^�;ť����"]h���Z.n�'6$�M�,y6���\���ߛ���c``\�ܘ
�it�l�_xϨ�j|w}�����V�m9������!���� ���8�ʢ���8;�VH|��)	�+�����y���p~(
v�`'Čo޼���/		����7ɣ	�v��y�R��S��HDNNUAm�pBfy�*C�VS�P��<0н/�~�tt� ��'� �j���>�������P���V�i)�>��W_�r9��ҏG�P)����j������X�uΌ��/��B���
���9a��	9n���#}v��Hv��ƳEz��h�L�:����5��jv���@� *�`\����PVHw�!@��H�,�@�(�O��r@k%��1--B*�2A$�1�;o�����Z�UP�!$n�ċ=����O|y-��.Ô�@2�Tr�Ҷ
B���h6����HZWm�;Bb;'zGG��G�M߉� ��|h��,p}�JҖ�����F2,�ar��ES�V���뚁�fec���[ˤ���`vo���Ct����4�q��5�r�b�kn^x�0�� e�g�~4�l�b����
�;�-Ə�Ǖ��z:\�ub5$�������CDA�J���ÅZ��[�oX�u�̟f�����J��5������O�H�%y!�WR���C���|��ŕ4K����P$�~U�_����Ѐ40�����AO	3TW��b`b��[]6��a��PQQ��������g�$T��u�"��M�����e�<X#����S�x{{Za��w1Qm&�/����kU]`"�)�w�h<H ��<�r�G���yaa
��5�/^@><���c�3 ��\�D(76L�1xȰ�u244<=?��wz����5:P:����i)O����Z�_߽LӉ�����3f�VV�~>Y�.�l�_z�I9�t���<S���bX�ύ���F�������J���L�,��(���T�*tz��8��ݏ���utt�m��$����}K�z �����QSScR��fq)(F�nANpܝ�SKe�32~9����j)��?����Y �Q����Mmچ�%r�3����,��@x���X�(x����ɩ>�[P����<ן�3
4>�v�V��Z����Ф㩰���!Ƒ!�������4� ����X�ht��ā��'$/�㍞:t� 1����0@@=v�4}u\V��6"!]ҥt(�!�}#�Hw��� --�]���t�4HK��<���_|�}Ξ=;�3׵;3� E���("x�����GIP�'ح��=o���}��>� T��(�T�	�U?�蚜��锾�)�;_:N��_���~�o��S�=Wt�7F};=u�?a0��-L���� ������-���@m H�J���ks�EXb�@)/�π/գk�Q�����X�>�y��5��4p�_z�[YI����<q��w�T�ݔ�D�5���I#���FFF�O�\>�4Ů`>��|�X=<�1��jV��~��)��~�Gn.����m ����$����>/f��w�����&��q� �8�N�`g7�� �{����=�K.1�{l y�N����C��|�&��;��Y�+tq�s2�[rr��b�{{{wu��-���p#�΢��B '����9 5O�m/,D �x�{��/mY-{�zb�h�������
����_j2~w���j�˱���&]���L����o`�
��{����H����d��W�@=><<�ӗo��'��G��J}��	��=�f��N�������//���S��j���wsv"���,z�q�hz|�S��`pbb \�z�M�H��E�ٶe�	�w���^ق���J���!F�?�g2�[�ãYj� m&pX�N�c�����������"&� ����HH���x��~̯|���#	�z9�
C�����_�7��2x<@��IIIu���^�Ù�4Q�H��ˁIKۛ�d����=%(���:�˅�-��i:7hI8�eý��(�(�����1�q6
��F]����<�߉�9L�U����}}y:󫪫{K��Շ�a���>@�;C8��I��!�Լ*BP��V�w��w�#���㋖����`��=�vGR� ���ޥ �D�W�'+��H��1Ʌ|wZl==y�Ix�cQJ��� ����,���Z��下L8a����lB�W��c��y��V!�7�!l�#	>}/�O�Xg�NƤU��$�*��=�_'~D�����V|�� ���q0�{v�ng(� ��,��2gE�����d� �öyd��Y���K������"
*V-�������@9$Mp�Wm1Csu��`%��jhb�i�/��t/8xx��RH9����`KW#b��^�����51�-��'@���N��qϻ�����V�)�G�t���P(T\J�M�3�U?�����XP^%hD�明���8}����m�����7:�JFcs�P�[ H���\p���$*u�!���&�n���t���t�3����<V:� �?��\�b�_H@H�����������װD E*����H�`�>>g����a[bai	��Y]U<�[&�v�����<bRS	���4����`4�,�M*�{c�0�-ֲ�n�0ٯa1�X^E�< �:^�DWUU%�|���7u���\_�\�������ӓ������Z�!n�بY
9�Ҵ��rXKL�� �gr~^2�Y�g^^���m^�
D� �f�_ ���lA�&)c���}D I�Y/b��:�#�����:1�-�_(?�4x|ږ�4�������,07���:��N��\�����v�����Elr2��\x82�6�/�<���D�@o��M �~���{2�$[7��`,0��y%�󝖋�D$��	��219�+*��Ec�LL ��l'p�D㍂�����7,S��+�Bx:Q'#�=?���oQQh-���SR ~�x̒u_�"����s4?2���E*�� ��o�(�D-.G��ٗ��#������B�I���0	� ���f�~�LIev�jP�"�����!��m��T56 �Z����$�q�����uk�{_�$ ڀ��m��a�� Z �襤*(��� ��� :����DaH/ݬ$���f��D
�����+<jjjRN�Q�� XX^�d`@���[h�#�����[YV������҆T�wD�����'�ݚ�N>>�T��� �P��Buu\ UUWwBK�M�>kk��T &4��O��H���`��kT��À���iEa���D��[������zo�6��ihs�JjV��
�ھ��Hn�j�ӹx� +��c�G��7kQ����}y�u���@&�[ڨ�ULw
�>x��#�C���ܼ<���vN 0P;����[[[�͜%�'l&9ykp=p�mt�Y�pg?��Y�t|�Υ�������6݀ԫ H,lu��I+�������~?���3 �Q ��_��~���l�����& E�
g(fL<Z����������� ,q�|�@����@n�f�`��䖔 ��r�t;>���qI�6oXހ�mzzd����2 A�6��住�������˿��?�|���T�E6ii{��+ |<{�n ��#����f�م~8��� �F�k�q����d� 2�Y$`�<�H��	>��h���P V���JŞ,��f���^"���S4)�F`�X�&�Z��C0�^��j��[0L�2��ю�Mv�[)���3-!2;��N��M����?�{��9<z���IO��4�����A�w�<�!��F�M�4�1xUs�P�8Z^���2�;�/�Q��GZ�X�M��L�����������lC�Ag��~�]��pސ���s�'<%���ο'g���20�Á���������F�I�j_�'��^i������MN��-Yn�G����?�-''G,�o�r'��mmh�Ԇ��6-Ɉ�k���cD�)�U��0r?,�P��[�%��v�ȏ�'y�y@����xxx Kk�h�F�����@��ڗ[�:�<%e�����[<�π2PJD
͕�&�5�D&�d������cJJ�@<�,�G�89F�ἂ,H�r8>��Z'u�ͭ�ﶫ-9N��`�%1��ٽ>(dx��\�gg�ʺo��7z��-�p�`���sB���%���x�cqi圩�pb����P(|�� 0�!""�@
�@�b�n�L�Ѫ��A�����A�!� ���t5(`uǔ�-�%�����Y�o�iO��H	�;/u���Db��s=�w �`�ziz�z�h��ę-vD�h�TvY��,I�DԤ�x�G���gƏ7ol�vh��sϩO.�����-�%z�G��o���ƹ

p��cf5��%e��X,��X'%�:�8�Q����Sڷ,��v4��\j�Ц0$�(��� 7?iuH�l�6�:�5�i�3�4��Ί�G��j�O��G,�����Ѣ�We�͈�6<�g�h,J�=	�6�i�̌��*N�H����"�#�4������&)�i��\^��1=�7',�yģ��g9�/�k��QHy�5A+�wC�=�>�խ-V��[�$�E��_%���a
�QSS�o���m�ۛP5=�<��vQ�٫�KJJB�"N�xr����!�C�=3����O���pW:23I�#bb�:E+�	[%$���fȘY2ϡ�/��CZl���Ėl7��Q����f�<��[�ju�u�ܖ ��q"K �t I���_�5W{{��~wԊL�:�3=0����q��
����C&U��&��#�`E���RFp�?`������/~�ߚS��꧃���Op}X��\�TfX/��󪬛�h�OK���6y߳�ȧ�)**֙O��E���ۦ03���8큩�緷�t������.�l�!�S��,�6\��B�]��Zq�U��n�ݏ���n0�K��0�[�	�@�6Z�����5�����N4Q6�>�P�x�Vד�P,J��:�`~'<YY�2����W�_5��}k����u�L�u-,��V��=9���n��U�@X6�u�E[����3�r=��D�Amw`�L�5�P��RË���@���ΑQQ`0\$�L��vu�����zW���b,~sztv�!/ۿ>III�c���۫�*��ܙ�"�<������[ޡNMM�11հz�eֱ��l<�UvF<sM���f\.K#�o�F.-��P�dĵ���MN���(VD��pMůj"}}x����� KjnU�P�Ϟh���nR�WV��8�����p����l�>r�m�^C�T�I����t7T�=b0DZ�'���PC]���� uY0�`V�]��d�J����#��t�.)��߭i�F0���b�~=~e��G�X*|\�&&��xV{o�)���o����4�yAF]�d���CC���$JA��6��jH�s�N���Xd�$?���=��1�9)�	���%�$�ֵ�`�W��+'���zB��|Ê�w���g�pREM[�Uq�p�O�m| 8��t�y��-��ԯ���y���I�T1�ϩ��}�)(��wv=L�t�~o�7	g���=P�
�S���7��01a\\Nt������c��	 ��yE'�?����(A ������\Ȱ�V��U���e��+<b'�;8�'0�%u�*���h��K�EWGߐ�E~]$Z�9�:E��K �у���( <I���mm��+�p�8������*�A�`� �:8�ZZXl�u�H ���G�Fr~�w�>w�K'�?�;�[X�/���t���o�Q�����ܥ���U�[E��w7eML�h��"����|i��`�z�Pcԇ�x5���>'9R�%�/�-�K��eG�M@OO�����Z�wor
ob�<�Ծ�&��P���K�0T�����ɉ2ʄ8W(�
�Y]-8�u����ͼ�?�V�6��Lu*k��K:������.u�_h(����z��L�$���Ó�x{�> f�,�uvMNb��	U�=ܐ�?�V����U�D��J"E���ӈ�I���/�:�%0�ދo4������cŗ��۞��� 1�/(����B�x��947��X��~���T�(ݕ�p��}� ۳ ���$\4���gj����A�Jb	'�"�@��+i�g��d���6r��_�fvv{���OH���q��(*/)
�[v�_�X�k_�!K+���w?������0�FV�n��6�y7�.�iaVF�ERE-1�܅vA�������{8}��=r1%%�:$����\t�s��p䪓���f� ���ޏ�y��ƗdD=\G�>������̙9�^Ȧ2͊�H� ��K�8%@N�7g���d�_==���t��f�}�z�}�s=01���-"��O�����xʱu��u�s�J�!l��9<�r��ү�r�t!,���,W�'="��2��!�S̠�Y��w��n�q鷧#��
������!�UŭPh7�on��6���yj5Tz�����_3�(L�.�Q���}F��Ԩ���P���_����K�M����#Q�ق��?>5y^3��`EP�T��^�o@~@����7�f�5!�V�Aۭh���e�*��wǾ��n�'��� ��\�tU�;{�eyu$Q���S��+t?҅0�ڽ��ٷ�����Z[�ՕsbRR���kDt�8��� >����ņ�l�ѱ1�o>=܂{Z���U�� `N�]NBM������*
�	���p��9�����2w�Pى����|�d�{}s)�'|��Js ����o��S����qx���@o�u�jcpg�V1,w���	n}y{{����Z�zyXYY��m��F~�%��3⩜�j�\���H���:f���`vv����^��¢ҡ*u;��!�K�4�M��ܨ��w�v'��lG䓛22��j��?���%H���B�����W����H`(C��69 ���N��Ů�4�p|�1T��aZ����=�IXS ;8���p���A��� *-����Σw	�g�������x���$%O��U�ƞu� �t��EL\UWA��C�Qv0�a��i�0�R^�*T���|�t��p��#��_|����ɐր��6����f�*7Z��!���W$ٯ�nj��=
�q@���/b�;�O�P"##�445���)�	��e~�4��0K��
�������ˎ�]�
;����n�M��^��
���u���%f������!�'�m����	҉�5�?+>;�\��ʓ���b�s"�d�ڙh�z"3j��K��=
FK���Dy��Ʃ�p?k��x����f�G?�X22$����㯨/����9Z�-���$�f'�e����X��j�px1c�ъ���B�"�ʨԐ�iܩ;7��Ņ�t��Q-�
ӡ;19,*�z�j���3X���'ˍK��|�((��S���"zΞ�������գ}h���Ԗ���a@X����E���u6�����������F~�{:�X�$%��}��S7�������k�����c��<C	�N:/�A(���=���ji�p��gS��/'e�X0"��� �u����1�{o���R3뵅��60����OK_k�2X���Mp\֔y%�3�|�[���^�5�,��A�%∭͑)�X|��=�]O�E_���ў�(l��ܹ��9?SL������0�����tL��0�\��L�5m?|�Pe2���v�7�(
�Y���1q���᭠򫩩������a ��=�����("0:Y��(��{�(FBC��\�0(��0<��h����p��q� 3w8���:��1q��`Q ���
���!F��&069����(Ɯl�)#'��uWZ�T���������FB�Hُ��-����ߟmʉ����1�SL�%;�3Ruw�s��X�ȵ"���M��K捿��r���w����\)Ӆ\��o��ïbù��|W��^6�쪰��=�<ZV������\,z���:'�Y� r����a)��� �M�|�p#��<�������#r��i�5h|�0��c��,K�Y��U:�% �\���M��࿌�	�QS���*7j����������LM�Mg�Be������O4 ���%EdTʗVF ko�$�UC|#@F�pLN��M�=O�y�p�d=���ڜ�+.��E.� �W}�%&x;�o�+�pc�6�)�T�D-��ncx�f�����-��c�K������^�b֩�)Z���I��❐�������Jޫ�(�y���Z=x���i6#ڟm%dho�|��,��+�!74LŔWVJ�ˣ����fgǠ�3��5��lG�p���y���RT߅�	���VQU�8(�޺�?sMς���l��8������0ē'���ڄ��c�����������}��߳����HZZ���b+�����*�duu� :�����M&N
��* ��Y�而u����PVFXI	��mzf��b�kb�4t޵��,Z^��>rHϷ�F�¾@a]��½��	 L��d�(%����� ����%�IN�6�	�|��+X��1����6S�`��hr!�v=�����	�\�� Vuy�9i%�V6s�qp�}�M��,��`~e���\�gd�����>�1�<�UWca����߃�-'�?j��|��#&p	�> �Gx�)V�𪅅E���Ǖ��Ф=7�]�����{:�R��I��l@^���,�lDyX`�-@����q�� o�&��	��� �7<<l�@�˗7\^��{��2�:��[����_V�Ӗkk�����D`e�큘�3���SPP�:�Z����w�2uKKK����
���VBUG���iM���~�� ��ć�_}+Aɴe��dxbh�2�Za������	?tDDD��V��j�*�g��ƹ!�@q��P�_�υ`�P�Ia�<��{"8_��'i�u�f{;���e��?pMD-����vܶF�}��Xo5�$�&]`����)z���y���eϞ�>����k�V��Q��=��)1K�����]y\�v[���W/�6�B��4�.�$r�����x�b�zsc�Q�ak�^�D0�\���YX�rr��x���7:K�W�n�7=w�#��{��q}��6i� H�r��#p����2}a��������[s��0��Cp��g�Uɐ�i���ce�r��h'
6F��ʲ�>ȥmD���R�	 g ���(dH�/���*\���˾�cKx�P����$�	�nѧ�n����hyS���8ZG�d(X��nV>���J���oM^��4:ޣiS0�cN���l@"%(}���K1� 	�U�=��J���{ׇ?	- ������/��A-�7����ˁ�}ʵSL��P��㱷��J�FH�6d��������5�{|����$	�����i��G��$ ����D{�1P��=����4z���kT�&ğ�e���јhrdT<<���S}}����3�Ᏻn�lk�I���xH&�v2Ix���Ő���r���t�b�ט/�f݁HfG.�ҡ�Ā�GP2�F����u�'��������lR��1�SU�&@�/���"�52���Lת��m�x)�}5T�/��#A0gm-.0��ƗإmuB�'�����Z��{}��|����R�ru�/0��!���cϥ=��u��ݯ/��"�T߿�g��+��~�۰_V	�O���	��T�B�J�F!��f�O_��[q��[{�v@�[<Pm�aL<��+{/u��p֞7����cSEP��5�,�,�X�V.ώ�љ'��=��	��7�G1�b/S`#�S%��h���-�g�E�9��7D6�\�~���Y���R��2a��-^���gX�]Y�,�nD�_@D� �y-/!��_M�y���s��� �e
 �m�ʟ?~����8��9�=~���;������Yy�nDr�s�S
?;i�|,
���0��kRctC��2v��}I���E!8�o+�F�!]���}�U��g��37Ov��F�ҽ�gbnd�T����+7-�ApbzF��j[T���^��"\lh�$%;�Iid2.����� ����J��0J���P�S����gec�B29��,��>�N7u2�f�]�;>E�`jWǏ����?�R�x�-��Y?��r���<9���J�s߰�o�/�b���}��o��`��
���z�pq͵��ܡѿ�$���	��_��\a�~ژ���n�Q��A�=-��Sဃ��4�T�:Ҷh��Z~bnʞ��?=��#91'`g�$C�/�ጸW�ǿ�!�<BO_K�?g��hPv�*�ˀg?��������q�L���Bi��	SO_ZQqsjk��7�8>.b�	��n���J;r�������&N�us��R��g��v�KJ�>jVώ�q+	���_�N��&��#��mi����}>��e�3~�˿����Nĵb	����h�':8�;������+���
�y��3=H�ao��l��	6��e�7��rnX�ho�V�{�����>	T[=8�ۇ�l��W�ױN�T������ͳ���%���ڳ�n��ڵWR2�F��\Fm%	�(�1��G<���:_sN��껇���=��a�a�����v,Უ�!f	�J~��m4$�Opw��� l�����Xx���L5�倛�3붜Q��(B�<����p�L^]�0�&��B��됕=��ECj���������u퐷�x���T���1���� :vp���o` �.�2���Ͻh�1�ٗ�P�&����c\n���jc&��g�g~/��׼����8F?D693�(�W[�Q�Rl�s�
]\w0�̋޳t�H�M,OLşM^�v�T�,$3i�����F���k:�.a"��no�-��pb���fG�2�*�� �/�Wv�𓹲ǅ���oy��\���y&J���{��+��O���I��l��U�n�ԥ)5�k���{,���HL��--9�1Fg~��sr��f��Chi�Crc��b����[j�ݒψ�VP�j�(-j՘�v:su����3��D	t�A���� ��!���/�ήr���J)�ht�f�;���V�k�=�������Tr��|���q��=S���n=�h&��?���S�x�&e����}���N�k�(6��U�<�q�P�J��`�1�::�4�(���65�S�^o�na+*�����]w��Z�$4��N=���ʆ54]#X��zta��Ͳ��ɧ��sN^��A�4�����yܱ�|�(��Ak��0:qh��1V���L_�)�5gm��Q̾� ���<�z셋1
��ڼH�0��$6e=͘��J.N.�/�?̗�[�Z^��\��$��*D�fQk	4[�3!��k�qIZ�6�� ��\��d������;Gֹ̚�^��˛���l{dfI{N�B�i����^��X���1сi����IYyр-���b���=?g\ֳ5T�2'�D�w��5���"�� V i}l0Xn�f0B��qNP�E��O�dwu{+)-=T����{���t���b��'�����Sb��;A����3��Rc�P��|P��bp0v2{�6�7����` �������B�q]�̗�Kb|��ċ�6"y:�y�d��L;��S7����OXXX�0�C�n\!h�e����ʔ���Q��G�!�����Sr���� �?Qq�憛�կ,��6_��>3�'�;9,`b���D���=^T
}V5~��+����
>�U2��/�$�6��ċYw� Z���[�ǿB2���!ɽ KW����u�I&&o�fJ|`��0���Ў����t�5��΋YON�������c��K$�ދǥ����|�Fxx/�d�P�;�덺���������S�S�j��{DD��sl���� 1�R��z�����Vr1QF����W�6�ߪ�}c8"��+��~	��,8���m|rpP�F�ތ�"����q$t)��k�8�G��SU�ܽ	S�Q�����m]���4\�O��&�ۏZ����bmO�I>��� ���4����b�����0�4R��G�}K�79�ǊZ�)�s|/7�K��v�!�3���i��Y̴2����`ƘHm�q�C���7���{y��SQfɽ�4��2_|�?����+s�����7/ՂW�En�z$�mm=&�����Ƶ��Oԫ\ok��WA�D����a�����S426�g5���)!���I�H�̡kSa���1���kcK��B�X@O<Q�Tԁ?�Lk;�����al�x�J��=��ωz��F�Z��G�7Skkҋ� 徻���d��0@x�d��XJ�����5�=�Մ�g*��[�ҿ𢐙��3��/R��s�Lkϗ�������U*�V_���ɨ*+C�sŗ/b5j��jFFfLuCU���ʵ�����&�4cB���=ZU�����œ
74�[�6�Z��Nk�g�u%��zx�@��\�Ӵy���̸(7�)�y�=�m��T�&^�-�*���e'�qq~2�.Ǜ���]8���Q�O��v�1�ta6�Mp!f|�Ј0��=v�~��9��S�Հ\lyͤ_����r��"�ܥ�\[�t���a�>jq�7lfb�W6V@>8��ޞ��&��_����s�Y�#�g��e0
>3��#*8o��ULc�϶LO�?��8��M������Kegt�)N�+ #�������_sm� ��x�6wy�3���;,�&�4��i2x�W���8�`�'5f}�$�S\�w���<q��L]�0T�)��VnE�9i�e��P%���c9�w����%M���E�1��[tN�쬳v��-�9�kBՏl%���L�?��g�Mv���o׆�k���06�Df���*	��jB�[v-����6���!'�-.�R��.�J�-�uPV�^�B�W�V�(<|׮�%C�}�
�{N^k=������l����{Ƌ�^�g�	t��M�<<��E�k�ޏ�2��cu����A`�������~�Zx�-o��`��+i$����F�T�ɳq�O#?�Ykv�O�I@��,�Q7ܝcDjN��I��јnt�3�W-�W���n'�m�u�� �|�-F��ߜ�=[��zIŪ��C���Ndiv�����o���U�B������+����<�_����T��-��1�l��Ƒ5�+�6�/� �1F��du��__���*�g�}o��2���A�$�Y^?jʰ���1g7ǔ�(T�/и�xH���ժL�徸ʸ'A�Ԅ
.��>y� ��>����?��V)�.9.�c$�8?=(F���px�؈nr2Զ�Q����QC�������a�I]�}��]�Rr����ل�:>m��G
����j�+�tM���?�S+���n	y���̺�d��J��A�ܽy�Q�^��D  pB�=5S�s%�ϩ-�_l]<~�(�K�=����A����S��8a{;4K�D�5+#Ht��qr��&���D�j����e�81:'W�Ȩ/�81����S)w^M��=�%e��tbgc��ԦHm�Y�^sVP���Q���"L�а9�7�Ez�w0���=�%���s��x|���2vbב���1.�&F�Ń�PQ�WY`&�Ĕ���X\6������~T�Ĩ>7�F���W�W�yE؈�h��`���nȩoQQ�v�Z�U"^��E�� ���e^{��;ۧ����J�$FZRI-���� �Ϣա��鞰N���rp��ڤ���7p��K��H�����5��%7ye�"�� ��bs�@׾|�ET:c3d\����!����� ���B=`���mx�ǖ���vi��d�vK���<w����Y�N.U�s}�d.�向,�%����DOں:�(.�K���gF+�Yq������'�j�ec�2''�w
8N.Ւ�6����n��_�.��פ��N����5TKtU��&�U���_'�v�`Fg�6^�%UR_�d4Ut��.>:�X���f�[�D�/+z(�t�k؊D���qh_�F����A��eq��I�<��A��N�����:��m|,�I�3
�2�i�x��z�>��!YV:����8��Qy^�E�ˇ"��_���\�7��망-��Z��d!Z��#���,oߠ;4e�d�`O��g*�@���p��S��f���T��J8>7� V�0)ϫL��@��O���%�H�T�����qq�����GR�"Ux��ϭ.�q��}|ښ&���>-f�#\�:��&��>7�����IQ�sS�kz�3'T��u�ח��]���}#�s ��Ҍ9��p�KC�m��M�?aˏ�;T�l���gjyb'\f==O^�ȌX�ឰ���63)�����YU��h�$�22�����4[WRnw� ��p��햜<�Rr��0Sg���;��0�|���;�����7���7\e<�"��ai��bK����r�!3�ң���lp��2����xT*��/�~��#k���f�j��iyݰ�3����lehI]]!��uҗMִ�eN���,��͔|�QF���c�>Vô4���P!���]�!���8��I��թv*��h���ISy�͉��h�s�222��cFvsk��x��خw1��^��-2��{EPU*�u"�����m�ȯ����?���b�T�k\��7�V��K>�'�Bu��Y��d�{n
xZ�� ��:���:e5_�wwѓbᱟ�VFT�:qU��yz(���PQpt\�� D�y�x�'�w�/��#t��!�%Mf��ך�NU��-�D�-�=5�����Ȏ{]le��
`���M��5R+�N�����L��ʒ?��|�����l��Д��2P���jib�/�r,go4�V�h��=��V�L�ϑb�lO2f��J��h�3��5_liZN#��5�k��WX�!�j��A���i�N-���R�r1|�T!L��"{�.-���Ι�:ڒj�i/	����*�ʞ��;����Ua�4[�A��x�eΒ4�&�GCy�)6��3nw�g�[�I��N#���~{�0Jl�K��f8\�Е���]��m�y,m�f8��G�O� *M�oܩë6У*0@p��]Ne�7P�B�ƓLe+n��L��o���5�%��&�r"��KmE}�l��-A���2sq�����XV�<C�r<ly�͂
�O����L<g�a�1��f���t<I�_���T0�'���mPپ�y(f�K����%iː$�n�0�h��:=%rfFȖ�3g���佨��pyϜI���q����M�R�E j1��Kl��FKfx=^A(�@���]3��kV�{`ϦA�ʑn�,~�ҒӇ���X�W�6*b1Ym���in�i�ﾏ���C��U����*J�8�^���EL�)fH7y����y�ZN7�0'�F��Ū�BD
T�n��|o[?-��9�?}��%�����v�ɯ/����r7 ���!,��|��q����p1�J��s��ںb�;Y��&���Yz���S�+����w"%��&���ּ���ww7g�U��挚tГ?��'��X_Jpܷ�M:Zt��L�!mj9��<cM����5.ᰣ�aƏ�W�!��^��L�`���z����؛J9
^���F�+U7�7K��TV؜*�2f9�@\Y�i:�7�{wZ{YޝV��`nyL�@���3�I�NvF�ާ�i7ƽw Zs����Br��*f�,8�������VX(�_@�H�En_�Mszog�G���PKYW���덳R/�8���م�%"�r` �v�y\�CS�32�~3��������G\�6cɡ��&��:�Yщ��vn&�(o���4Ä�n��ϯ�2�E�;�j�ҳ4�:o�23e�LO^�q�x��9ds�(z��9#�"��,U�B]�CWұ�������Y�?ϏG(Sń}��a���6���-������U&���2�yˎ�E�Yr#h|!t��1s�
��ce�~p1F�{[h�Xi)��ȼb"�Z�?g�g��Ո|�;(�"!��W3�w`"�����m�j�)*�p��v032S��@������8�����\�2M���ɶ`wjZ����0ԩ�88JO��K���6�c�*�H�/e���~��G�8�JKI��޿�����!~k��q$Zl����W�Ӓ��EPIIp�eg]]k��'3���/iF��DF5!��B���c���/�/"�6�9v��Ŧ��~L��Сm%[_Z
^
L=�_/��;~�;���j�[[�Ե�r�7J��We���`5��n��K����~�@'k����f)P��������J�n�|0��b��� ���W���\C�K����il�A�����ٙ��ۺ���Ӛ�*�$��Z��Ԩ�˅%B6+����RvC�4����T435��4ι,έ�v-q������ZxǞKc"�r[(_��Ffs1�6�Uy�+����tn�q�ʍj{�&$�m �d�XL� �'���@e�N���G�G��Г�h���ޕ ���35ޱ�~Mmj8x��p�1��urKE��Ăweɕ�D+lG>�kؙ��d��u��Pc+[��R�����X>����&J���ҟ���Ӛ$O��r��ƒzo\���+�I�w�0��
_�s���I�������]��4Qq���{�vi��VQ��0�����Qk��U��p����c��no˺XM��#7�Zۢ�`�d�~�℀0ʆtm^��xG3*����
M��{Mփ�a���bY������7�{�䢐�G/�Z۞ɷ���Z/Y1�eg3��#+3���@���fQ��K���Y�2���s�&�e��$=o�=`�_��kPNS 9ѧcZ�Jb�%Ol[�ޕ�Q���ڔ���#y��E8Cw@��$"0�~V�R6i{UP���翝ԛ�ݹ/#h��GB>�`���8�{<���B�����G��z���ΎђU⊂l�5��#�(��"��׻���?1��S1+��.�����HH�*wY�D韜\Vfm���82tuX��b�T�Xk��g�	�(��Vhӧ�Թ2�1$�*�8J'�qs�ϓ�#^�o�&�l�jb�1��|*t{u�kUَ ��(����N�pR��T٪�;)���BM��N(C����$0�z��C��z�C�у!ԛ�au�77�-:`kأ�$0VuG���AR�э����|6=P�M�s�BH�Mlr࡞�����o=��ޜ[b�[������nwU�nu���&�`�i��""4�Z����+/m��ܜ>�~F;��/jű<\(��L�)�{isf
�FNf�ۭ��i�=\�%�Pz�Ծqz�ϋg��P�S]Fks e�m���O�*��T9:��s�������a����s��.+�����K���W���
��RSs�j_���ywO�\�8`C�����]�ӡ���0HH���&��+Yß��]�"�w����I�謵�����c���f+6OJӻ��"�	�T�|X�Ng����9s�Y.����n�`x�4��g4]B�%u5��Gzj�2�!��7Z�k+JK�|���e<�^d��de�{��'�49z�7UĦ��(�a��1[ƙiF	�&MX�s�^/�H"�x���]B�]<).L� ��@�`���Ny�:_�]2Je8���_1���;��Zē�b��Q� ��]S�4{�V��r>����R���m��ˀu|�DB���ͣ?������}:Y���>�Ih �e`d�;[��*:w��x$�)����Y"^���e�Y264�ylP���Ӥw�8v�,��o�\��V`�Q����L��q��^�0;�P78D5f%w�U���yN^!�� ��|Z�;Z�D����B�&�ˎ�-L7�nr�W�2I���b|TB������}����<�_oucqtt� ���V"W���\�٘�"8���8�J���9��z������*p-y�U�.��?zz,�4��F]�՚n�C��&��<A�zY�� m�>�#4X��j`p� H �8C���ÿ�'�zF�Y	HH'n��aV��������o ��y½I6Ɇ�ٍmsc�ƶm�bgc۶m۶m���_�W��Tݙ�QO���9gzg<s�/��O/�;J>�z�q'���|�3$��R}�B�B�V9�SR�m ��m����䴃�1�~�Bk�!''�?����e���{$��	���83�!'��lx��l� 4E��@FUa�c���Ig:���x�J��A-�}6NY���
3*����B�ew�(�b�p��2���G�Y����%y :6>`������l���d��*Y�Ȼ��j�� U�v��L�M��x���o�2�t�i�e�0k�8��I�cɜĦ�%��$~��]��
Ƶ����d�A�a6DOxH���/N.���	��CZSV��;$nbpX2�&��&�.�)ٚ��*�h�jB�S_��=��6>AM]]g��D�ظԨ,2$u��SSy8��:޶���o�Ƽ���?9�s*�<�̵IEc٢A!Tf $���G� ��Q"��
k7�$�a�!�6oM�6{*qo[��ֱt����Gu���dQ�ݛ���YK(��&�/A�8Q8X�&d �А�>g<�J��t����<2������H� �U]2��kʎb�P�+lq`#���&+;^(�^�s��.7��|1���+�:�th���|�}7h��Yh���/��`Op6�4���{l���k[% �!F{]mq�$�tx�Ȃ�F�A �$߾<�OKP+�y��|����K�k�<	0"�V�8�Z�̊����L�w>���Hc5����m����*�Bv�����������0��"�h���g���gE�WH@%
�[?!mk�L�s'�NR�ہ�hP#�Xx{RkT�yu���!J����x2x�0� 2�>)K�3�u�3R�֗��@`�,ˡR�Lj�\������6!��w}���� �TJ��)�Կ�a0qo��H��* ��j��ܼ`b�@d�7ffV�Ѱ{�C�͙Rd����� �$u�ꊣ�Z5G��IC&9��;�� �	a~�����ǒG'�{+V�p\�|gW;H�u��!2H�T���15�� �d _�}�T���'��|�T�'t%�E�{Z-t�����K6��+�q��q\�{M5d�AB;@F5�F��e��'�� ��/���WI9� �x�M�Z��x{݄]up��
����2sc�d��8�y��I�V�rm(�s5������f�D�Q���#���Oc`���[�Q<8N��Z��j�U�f�W� DlN���F��Ոb	�)֠�� HY��Y���?
bj�r�/xʇ��P�Y*O@�,2CO�h�.!nɑQ�]���Ak~�ٙ�3�)4�;�V�xET!݀�b��b���c�Ydɔ�9��T�-B�G�))��:���ݬ���ܴ�I0	 Q��f�L�����3�b�@�iC�̤��T[�X��4&�,[$�u	�!Vr�(.	N����(-�������Z���z!�yA_�	ʞΰ�����m7S�_�Y�UMT�r�y�%ye�s�L9Ʊ�}�Fhh������]��Y�y�93T�_������K(f�D�R�KfRnv����ﬅ(>��v�����������}�����k='M���"�ʈ��8e�����{3��?�s�"��E�䊅�f�s܃�5:ҀZ*e�D��P;����q�s����K�i�Wl>��i�2�/��pA��{�2z��<�Ef]��>Ӣ�]y�ۼ�'����+��e��ߌ�:�fgo?�ml�S؟ݛ�4�)�~w�8c@>]�J���;κ)���:/�WW� b��uʡ��T{_�����Be��G���9jN�[��oȨ*�C�ĺ��;�7!������G�k���o���#�(��l�D(g̫��2�K�F(qy�L�!�|)�yU��ɤaB���c�߳�HKpCHP����:.�)I�tw��՗��s�g�$��[ �W-�o�=�&MާWc� �QIAq�:�e&5�+6��9R�B�Xz3�3�RTn�k%����tB�ԥ��U	��bs"�����5�)y4-C^
J\�s"U���a��"����3T��cGl)�0%���ݾ�S˂�no/Ɉ�J�*)I_+d�U�㶒3��f=K�[�?�/uz+)< J��)q��M�Ԃŧ]]��e��nſ�2AnXJJğ]�υOHA���d*H���,AL���5�@��$�b'G��ye�~щ��oH��2W�F�0�F�Aߞܞ$��m��7+�=��7������+4���'	%��zs-�CV5����pqV��I���^y?�>�ҍ����mģI��bv~�$�g���1?M	�viAe�nĒ�q�<o�5Z��/4��^�|���v�i�t��5���''�p�����P&����My
��ǕK�������;��b84՟�����:<���2�rgN��Ob�w.SPm�V(�:7 Q�k��;�'��cο�&��y��g����ߖ|����'��!�����
gA�6�����L���N��4b��)E��Ў��ޙ:��k~��� >:b���1u>tp�g<���b���65����D�E���.i^��V5
Y�Mpe�"w�Z������Vo2dy��L���1k�;*��Ɂ��|3Z�4�@��"G2��\X?���%>�D����}{��A��>|ơ�X��x����-���&P��-9.��'�&��?�
m �%`��0����|{x�O�F�k{���Ǝ��MCf�?�y��C�k=�,�78��K���gw���۾u�}��.�j���R���������Z�6�`|�b�J���;)����U����6W�쎷$`i�$O؆�GQ��F���\�Y��ށ):\��e��ʷt���@M�/�9�<3��A�\p\�(�8?����m���ɑ�f���S�0a�b`>����f��K}=H�eϳ���@!��k�l|Ki)�Nr�������_�1JĠ3.TY�u��&~?�թ%�׀�s�D��~~M%�[?���_X'�+�n�U�xh�]���s�ל8sHB�%$,�N	�U�4A�	��
�CA�].T�Y�:W4�� �{��w*�#Ȟ�"\�Q��k��tHM��q$��O,,N~�R��z#��BJ��vyq!k�f_^^^(`��a���/&K�/m]er]���H���c��C��3'�y�9�h�y�é�,��h�^�[��GS|᱄y`��c	�.dM�P4
��H-���G1�xV��9�"\�%�QY�w w�\�93C��������퍯P(�w<�&Y��s�\�R�V���f�ɕ"�͵I�?�:.Bڏ� ��Y%���O����)�;�G777�&���Q�諦�v�؉�l�6�)�Zx6�	
��V���\�vYtM�4�͓�����2�煌��b�j=��y�B3�N����D�U���8R7Og@����L���T��E�����37�v�7Q���X�m٨�R�/''f�+��rW�V�d��5���gV0V��>0r<����>ҽ�Γ3+�-3�4ѡ6 �P��e��Xc�/魦~:�T` ��e���A�0�_S�[T���h-��P#��mh���)����5:F^v d}Sǭj`I����n��Ɖ�ssRt������pw��y��j��ײ\�nS�98[�A醻8�I��"���qSf����Τc��K�;���r�D8��[V����j���p��6�fKC�Zf�Og��RpZ��m����7��orޏ�ܨ�t��c���*� �'S'��kxc8�
�:A&�!Vuj��bV,���Y]��b��,���jtlY�� ��y��� �t��M���./ǅ�22���W�gw�|!\@|�RD#U��1hgz��7��,������vH*.�0]�=�ii�q��H�����c$���vX���MȎ�J�W�Rժ��gC(`��� 7�m �;��ٓH(Q�;��.Y�Ƀ=�^(�[�Oh�/[5ؠ�_�G�XY�&�5XG}����poA~e����\�ޞ��vĄ	��U�Ab��Yp�#cC�ũS�߄�i������l���������?%?�x+UN�g���B�]�z`Ìs�)R��؉�w�xM��'Zq:P���=���EAQ��,��犉0L$ԝ�/��0#q���"R�zha��X2�8�\�3�Ռ���0��`6��	9@�U[F~ �c����c�Q���5�Ә��ί��	�1�K����wQ�0h�� bp��� �L����OP/�d��q�񺃑�lGSU����aR�,��V`��|��=
Q�F��C�|���<w{�CYY?���`X��puuuُW^����s���L�����v�����E#����*�ا���.��z߆M��瀯e!g� �I��<���$	��;�Q�ȗ����<=� s]<V�����i�6�g�'{�����G�)n��{��N���^5P����O��Ԫmb>��<Ֆ}9��yj0tDJ	ʽR�= e4��x�r^�㔾>��"<��,�(:��<��g(�|D���)y��+�����3a�k���k�E��
�G*?oUi�F6�?T��ٻvԭ�h��Xu�P:@ٛ���,%V~nW�����Į��A<B{�M��,B��/N�Yq���u�=A3B�L��O��mKK!��r�*-OX]� A~��z��E�F�N(��j�}�"�.N}��ޠ���OϾL�&d��� �{7���Vx�n��U!���ǿ��yxx�����
��χ<](��a�-?Û�@��"������=?�]s�uO��U-�l,� �޾�!�ScmU]��aT�б���&ņ��c�6��'�*r}��i��b����f�bf��!��9�W�O�|ۥ��	jf�d9�<=d9g���`bP��p� +�NG����z�ʖV�h��@Q��2���g)R�b��$匽h���~T@���ؗ*RN�:"���BiI�H9����z9��x��(�/���P�v#���*/�(?�ѳ2�E<#��E����3�''bb��V%�����j;�9�נ9��IG;����e�0�ժ�@���+��@�?��Z���#O�����̗(�+��p~8[~��ܝ�D%^<`���y΋~�:Ȓ��ڐ���e���{�S"�-}���v�؉W�6\�uO�����������m�MM�s�Ţ��!�G�+��*4��t2���߱�ڵ��J��xy3�7��h�V��!�zI}��[���˙�ˇN���X���_���$�Y� ��X��]JQ.�Wkn�M�7 ���#A:�2�ۑ��cdP�����y%���gg}�5�Y�締�~�O��ˁ*���gMO��t: BW�^%��i�,'h�-�*Åw���lؐn�T���ծ4�#�f�{Q���N�H[l�5��mt��QQ�8&��W-5A�����|��	ps5�F	V3��_�����Ŋ�#sҏ��.7��dx_�O�k|EmY?��D�eA���'8�s��VN��~ �#(����7��U����uFF�c����0���Pd���i8����rN���:=}���6�|�w�D�����g}XL8.�k�mj`	|�����$����o�l�+p�8��Ƶ�Y��A*�wl�\�����W��h���]�$D�/m��7o��J��+�����~״BH�����b������ݰ6�ê���J�i�H]PP���q�Y��38�8��h,k�L��]Rni���q;Wߵ8�V	$A�t�`��%g�X!
k�;R@O�Ii2�����(67rx�`�ONN��t͵�A
Fg=l�$)�":��輵��01�s�bq0�Z��%렺�����ZنC2&-4����m��/bŅdrhc|�1�q��}���"�ͧ��۴W�hԠu�.��j���?؅H�*�/@���ʇ<a����0%�(�ơ�$�x���y�6t=���Up?`��L�0!����`|{qO�'E�c�� �@��ذ�����U�Ki�M����l|�0�a�P���:)��i6m���24�a 6s��RO.���]�ge��G%Iz.�D5>CIViB�2�x��׮Iϣqpv�MII^A��lt���BT� ����-!0�uOeVJ0/�G(���#l���j)�Y��'�(F�|��:5�s X�}����L��3D�*�6�K�$�S`ƺ�o�HP�Z�Rx8����]s�����+M�*��96괎m�_�F@Q]�b�����+=^XF�ח剴��ؽ�Z�8��'��+/�����<�"��;�J�]�Ҫ|��bˁ��(��)Y8���\�_�Qml����_9�I���Q�� ��!��[���
�,]��4���I�II�H!d;t��s>B�Dx �\��y�85?�'�����S��}���E$��92����Q�_]��ٙ0��2 �DXP$ir���^�9�[d������r� �9�?T�]J�g��;|����ָ(:P����>s��B�l�ae؝�Jƥ�E��8S -2W:��4/��䕶l��VX�3���E'E�tfP�YP ���9y��i��{|�2��{@3"O5Hh�H��s� Pa���?CEGv|:�IIj0��n��A5Ho[�FpN�٩z7��S�����u�n+�ȞuW�ᦕ�Qi�)EVd�5��u����^[�ᦓ�-��bS"�&wJ���Ⲕ-=!!
j�ꉘ��
(�����g��01K�
K{8�Bwȓq11��>vʷ�%dh�EC%ʀ�]�?�L�s慇������ IY]#��|w�\��5��>?�	��Q���?��*G_I)~G����ޟ."��qm���4�q�y��F��-��Kԡ�9��z���E�m�g�k{9)es�X+�x`��@u8�]Q\!�7`gq�����b���+��3�kbpX�]�j����tK8~���U������9m�W,���?Ӧ���]��͙{�AA �}=[�][Ǉ�)K��+��kb��oƀ��6� �ÕX������`��I���܉Wv�� t�9W��9PҘ��`��ڂ���+C����b^�WŰ�`��"*"�c�}ϔr�U�|p��k_�ʔ���KJ�
a2gVq:D_n�lRg^�}= ��0�	9=����T�~vxj�i7|��8���O�8I�!a�<��e�t���	��[k�@�+6Ó����ɕ�R�) ���@�5��+*���Ϋ��O�hh~u��ǽ��߹�a�Ml����������k����$�����4�J��/��W�a'<f�5(�������U��
����o<�@����p����5 �塓�N��������m�9::&�Z000�bc���1qݎMEt��@�}N#�q�Dm��
z�Cz}n�`��;�N�~xx`�������x�O�ty=o��h-S̂tt��͍��������a-��͵!6#q���1��PPJ�yr�u�z�=��'*�=�F���=���/ �@B�|P1����u��r�Ɠ��k����ލ�m��X�X�swgCD��W �l[��,�$���;��0Yh�	�P�� �+�ν�P��AfYdD�z[R���w����Dĥ����D8s�����H���}u{���tF��ӿ�q��?��XYc�����ƣ�AԵ�~/A*B��ڨ��~H��ۙ�����Vv��	-1�1��y�;v�W؇�_6ަ���[�렍�m�Yq���c��|`]h-:�F�Y\�ӳ�z.���oOlޤ�!j�.\4m��_��]<�$�/���w���К�EY\��ݿ��`K�Wb���J�����5_��>�[�y�S%?4tN��O�'�rl��wȁ�I��z��t��>�
���m�CMA���D�D�0�������[�֝�U��=}\o?^m~�G-=�α���VN��zg`5 %%�gfg���[�;{u�nRu9-oĪ�Æ���`/<�a�~��?�"�u��x��x�B�i�Bw8����L�����"ؚ|�Z��X��o1�$���cy�G��B�)&Y���-"X�c ���:����G_�����v���u��7��j~0-�I�(��͙�i+��x�}l4d�� t�
~m�_/�UoZr��n�)*��gG��WH��?8@1p`�&q�Z���8#���\��&AO��nX%w:xL�� XH�.���V���!i��_���YSپpL5��������џH�T,���b���W������n�����B�|�|l�X�'�ru��#W �"-;<�+ƀ*ޘ����x*P��V���,��trw� P2�h�����+p�__�sd�4x P��V��q�֣�L��R^�Ύ}x���`o�P��e�%Ny5"������<�pm;�1dT|�8�E�ߝY���C�*o�7�+^�(�b�7[j��=98rbȘ[ �lh���k��]Mi�%7�j�D���*�Ҹ�x&���h`@%^��}S�:����ٟ�����B�9lz�	TE*Y0.{:{�6A�ؔOB�6�(�k�8���BY����UL��9�N���W����s���������!!!.7ä����`M!7��F��^�7ؓn�:e$x�P����o<��WB����&��(������w�un �����ȩў�A w���K�����~�g�(���z WTRRPVv*xsV��0�V�H�?�s/�@/ׯ�F�W弊�0�s��!Gs����t�(����,��C�2�̨T�oy%u8�gs-��!��c��T�0�}~)�u{��H���**�ͷ\>�ە������`�M�^�]\;���*RH��J�p��W�@�"��޵V D<)L:�ј�b�5 �KiHO[
���Џͽ~�&_�D4����}k��i�K�`�1��C��[s�JDj�<ؠ�]��'�΍�֠c�;���P�	�=C¤��)3����%z���HGL���n�C�T���L��@��dzlM~�������TP��E&_|���n���dv�)�� �d$���ڱ.jr�_ ��*�C��Q�W$��w����#OגKي�q� y�����r�Ke���q�)��V`�X�a��R)G�J6�1�C�	`ߣ��4h0��}��2y�3a8����P<h�·���Ʉ�i[��I�m�5$ឬ�$�hQ��GH�����P��mIۣ��cC޼�wm��	��
��x(���Y���X�\b���c�rֈ�D�'y?񾒷H�"ab��,]]�457�����F�Ǐ(���_i`�keRW����J;�ʰ��������p:{H��wn��a����~4( ��}��$�ibf5��z�{�$�Ȑ�X�:#_�������X��}�
�����퐷w��`�ZA�F#x�P�єaw��짓F��SZ3#	�z��9m�$��ѿ�*���S�f�T��6w��H�jѡdF�����B�y�ܞ�{8iA�g��L\�ţv�����D��A������f�n�q�����g��j�3ħ�Q�1w�c�� �����7d�x"($�I�E�����Vce��`��k�`��_w1|?� 0���ČH�ĸT��y`&[�h��OS\/;�	ck=w����4AB�\<S=cLa�Z�;wiMG>�2���Qe��Jٹ�+�Q�R�L/So�!����L�.y�����7�������{q	���R�\�6�h%*���z�h[G����B�Ky�e�2��~�ks���4{�����ʬ[$P��Њ$M} $g&�p�^�-��K��!��s�os��!��ʗ�dgu4���9��p�Ŵ�z��Y	['����t7\\�\k<�텓�/F���]�`���(An}#����tW�f:�B�ū/���v������G>g��q�����kL�qq7|ƌ�&<>]7B�5eL�xY���
^����XR30��%sߏ����0�8��f�tR�A�dNV�ۧ��JhKy��z>og��R-��N�C���7��uͽ4�����y30�� ���-omVq�_��v0qi�6�v�r2?�GÇ��Ie2$�!ɔ���UO(���ܻ�e��w�99dp�W��SL�
�����]0m�ug^�'�T*H�_��Q�@���r�ㄵ�, |�C�)`\p]e����ZQ�A����]���_ĊJJ_�����	�����)�~(���iw.+���u%N?q=��G��D�ŷ��iieVO���l��,^�P��4ٶ��R��h�,]��G��������k���ܲ����^-4�hЮ���-m')��*�������)2�.�u�W
�`�^f˙#J�S҄���*Ϛ��*9_��w����2xI`c����ӗZv�4kf���`���hRi�촦g
��ԨlY��=����Uk�Z�	W�ҫ���8�	@�rs֮\~��ٳ�"�,�z���7ؤ�(=�r�%����N��]����ً�rs�:O\,~����v%�ɞ Ĺ���vk�'��?���r�k~�Q0{�o��㿕[(��ݱ��ǖ^�S���hW,�X�=�H�L�{w��*�Mv{ZK�r 4�:���\����}�t�gyAG��کL��X�Q:.+	S���Zy{���D��i�i=��`�e
,�� G��{VEE�m�Hv�Xq��`$l��H։�����I�����Y�����ŀI'��٣�E�:�Ӏ�����4a�����\�'�q�,z��aZ+&8T	�=E��(0͒	����ҝ��j�A"t��t��	>���i_2f�Px,���sQ��\A�5�B��U��/Q�{��L�l�ܾq�#��YMs"K�Z9XԨ�(R� Wܺi�x���Ԕ�f#��@����%���/'��v~MW*�gP�7[�du� �B#p�tUkq�����ӓ�E�-�u� �<�I����"wꄚ���wH�o�������-H�=���6���˭�~��KX�YC�Әs�-���L�����������ґ�ys����ќ�zi��� �6j��P�*��Z�^��o#�K�}j<��;�x>,
=!��\M���FA�[�Z��ʔ�ǿ]��a�[����� t6ˁ�9��c�����[����Zk4�� �诋߈((`��eco�WG�����G|%��Uf�?�3�Le�)�` N�j�H̲�[���;=�����H�L�P�5�x��H	��3G�u	I	�c���IǢ/���Tm��	��ci$X��YK眜�v�EXʫS_�K���~�iv��LY�>u����3������s]��|���|�51�]8�b31��m��޲-�=�U��<�!c
5�O$��7ۣ�1��G��:�� 4\Q�w�' 7�"��ml���n]�;3_�B��[�4��M��6�sи�ɩ�OYz�'2Kx��Ơum˦���D���W��a�&n&����I�"-�3>]ͯ1l�ZQ[T��;3s���@�ǲ_��ٞOЖ2�X瘌�x�v�텢�,6���Cl&�3]S�{KQ��o�B��\������1�O�B�̘��i�úF�r�[S㐄z��q�*jj�)gbr�r��}@2����-wrҐZ�c�ȶr�;zE�}`>�52�������&��ЊX1@�㣢���_�V,b�SΨP�_��_���S�FfG+l9sUJ~s*�n�dD5�_ӛ�q���)� �x1=3������)G:��i�s`9�2�\��a�TD0��L��13�B_�ݔ�����n#!ێ�~a>�������U����<�,�ب_��Ul1T�-e��LjC̍����ioK�߶��b�H%���3���*yi PR4�����`tP�H����Y�nz☙�����@ǰ�x3L�N�����bͿXY�QNKiF�M��3:9꘮2Dݩ�f|#=3k/+?؏.��,[a5wz��Q�'s�
�j\��A�����]JUR;q�ą�6�����\��v6O��v�Ygى:==u�P&���A�hg�CS�}u�&%3%!McG�Y0G�p�Q=�S���<)� *���-3��~�d����#���S@\�i~J�v�pہ�Œ<9B����d0�k��H>�����%E���MSM�4���z[��|�#�(�����[Z�F�"�Lfp�|<���T��Ύ���_y&,W�pqÊ�����t.7�M�XZ�p��$���}�t�$�����0?�u�f��~��F������]W�g��a��mFoO�QW��"o��n߾}�_�U^o���U�ׇ�O���9�u�7	b6�q�S�O/̴����*�Oߜ�w/L+����ڀ�j��?���)��U�)�ů/Z/���q�����Xg999���/U���z���Ӳv������?ޑ�C�K�C9� Q4���5x/-7o�8����&�?Mm5�4�9��)��z���$��hG��lC����Uuue7�}���o}sљ��D��	���BN��Tⅳ����b0s��T$��d}����.P��gB�Ff�
�$�
H�?bXhnp	i��D��?�r�</z=vਫw�eKu��c4 �z22�V2�#�#Q���n��^C� ��s�|��m��,z���˞&��Z�Z~��� ��-O���q����8���h���{´?B�~4Y�o�w�m��8/�?�����{\S��,����݈�W]T�S�{�8�:�$%������=��B�Xr&O�"�;�S+Y�K���;��	�6�xw�rq0�)�V��w'���e!�6sV���|����P=����13�98Rґd�a�!����/n.z&��>��
q��`c__�U��*��ڠb;R}�����5z֛�֫�e�q	}Ǫ���J;�<��i-=�ʾ��m�{^��v&�{qk�TQ�[�,�x�	���Q�)paC4G�٦nMy�1��]ć������􀻞���]�P��f�p=]��>��R�Z]�x>?�N��u�N��sc��4�\�P���dq!ۼ��o���?�
�'��5���Y�*V�K{,��-f��A,��;���V�=�FIQn�B_/g3�z&������s3\��Q�6�A���r����+���U��Ҡ+!�������!^�
�?
����_E�P�vbO�v���V�p�g�$�lRXɺ����T�C@�����Р��M�A{�V�a-A�K�o�v�^J��&��l'f �$CF�zN�a��t7���p�3��G�׏'.����T&���{+<VR���Ʉ���J�]WB�cp��+W���B�E��칽�G����᧝ÓZ ��Y��p�Y��C2�p��/�r�D_�ي!I�����ǈ^�v�z^y�� E �r~I"�(�d�O�:��!��a.L5wpD�d�z��m�N�?aC���;�+�gex�7�ݳ�;����]9`��j~ˎ�c����СO�6h�J�M��:,:��S��ζ�~�w|a�mDā�z���J���¯������7��������惥���	�������kh����a���%d�^���tm\���Ҁ@���E�:�9���ßԩ$�-i)q ��������JĒ�tfJ�.=�r�XX-x��\>���~���C�uf��p��Wd@�5-��ԅ�"�|������ �{����ݽQ�q�z_2�t��5��`�n�O����rQ�@�ƹ�����'�þ�2��HTF�6e��M@��㳰E�(|�9p^ԯ�8e9�&cY��ѤK��$��,�eH�)�;��D>��BK+L�u����xq��G�e�Ȋ�Be��	��4�*�hf���x7��e�7��>Z��'@�_�Zj"���%bI��g'D��;kѪ��;�8�hV��	,�k�oo�j͐�3�w�a���@H�p��j�4�i�w�F��n��n�X��0�M��#��ŴNMQ��yq���H~�����P��|��b�頔�*�x;{�b�
��ln_�w͸z��	Ά�#Q�`]&w>'�����c�Ϲrg4Ȑ�|����U��yz�
�R4F�ё�j�t�����'ND`��:_s��b�+ED��ҫ�[�����h��ئL�텭6�.E�l��-{OG�C-g
�+��!_*D����G�W�7�������/Z�6���?��k������x�Y��g���L\L�Z%2D���*�������~!��]�˪/�fb���9��	��#�	~:�ӣL�\�?]jiii��O�͚#|f��N ܃��k�R	-">��N\r�Ѱ���z�ԛ�K�r0����рH�A���fّ��u�P��|�\�,�8��P�^��r�?�3٥ޫ�~���B%��p�>�;l���hJN�7~x|o{�7���-P̨	\	hhO���-R�HA��H<D��y����N��z+<�g��m��=���Y^����k�a%
�
\�ܕG'�}m���pA�_���22�9W��|%���L���=Z�˲��=�!����;<�Ma'���b�⟨����D�k�)!2����+�,�}L|� �ԙ�� ���|�����?�c����%�uCz�ܟ.���vOLH�mv�7Xt���Zl0����:�̌ʗH�;�+���e������4ȫ7�@����aH���l�ʘ;|��Ȟsv���+�Ŷ(`��:`WhO�!~�sss����c���J=�Q"�}:Cs�r�V¨�--��E�0)u�S��5�oj�+c�]~G�D�ѹ�#�T�y
\����c���v̱�uH��N{cb�|�;�۞���q�x��<)&K�p\���}�J�>lE���tNƆ�;LJ.��+%b�0Zس��q��� �F��󔯒m3U��}t�X���z��hZ{�V�����}���29!GOT��+"Q��С��#�]:�k�Z>�A�.}�@Ʋ���u�����;��S�s���V��s�<�i%�1�M���I�%⎑\��y-Z�O��*8ئ�*}�1�E��}QG�'V�VT�&�\�>Z|���W�n�RS�Y�:�M������4AAq}���Ɉ7�REo.��6��m�<+.N�Z��ĕ*Վ�zl��4U��]�A��P��7���v��\���o�%��?���֖��Me.�Y�?{�������f�#T�	��`_s�+;�s��(��1&i ����a�/'��j�>���أ�V,�g���C��Lds��L���[�:Iyr8��N���ZY�ʝ0H��.�ryޯC?>*�@���@�N�Hۛܽg�*����*�;�C��Z�9�7�7����?N�!_�d�ށ��}'�ԕgmS&5�]֋���ׇs�6z��cR*����E�V'ꯃ5EEşLsE4n���YH]�Xjq��W[
ƀ
@��P��7�Ϲ���@!`��.L�>Ԅ�G@Ų�NM�����,�c8��~q���a~~~0E�U^򻛛�8r�*�n�dFhI�{V�(m�gb��-��Ɲ��6.b���#$k��=�r|%w�������9�bzE(�On�t�hxd���M����"P���2\�m���sy
r��:���^/Ng��a9A0W����t_:��m�+�C	HȺ �+�q$1GN��)�,���}3\n����7#5j̿�zpO.�-)�1��"����q�A{��k�4�<nA���y��h�uU�ʨ�TBO��M�
�<龧�ǽ�^�h?�9�;�V�����
س�z��̘�K���}��[�eˈ�J�N�&�d���*�7T#B�7��l�|�X����@����W�W4���Ŝ#݁H��tF|
��Y��8u���Z�P����'��׳a����H���륜���़7��A� ��Gk�x�Qki]��U<|�/�oNCF*����;�@8��f�0����j�}���$6[���o��S33z�GVVVI��_��&y^�	���Ι��L��x�p���aP�$P���dum����QW��4���Ҷ)68)��lw2u��A��?@01۷���_ƘKae�#'$"��*6��,I�hJ���@xQ���z�V��w��=��Ð��e5\z�dK��k��ʴ���l��۶����ƙS���"�:�G�'ӧ� �\��<��� 
�r�:Xmd����������̖�E�Uei��?�z�&�����0�������ՇY�����R����X�}�5������,ߩ�ӱP	��T��:��+��	������;�~�mOU��y��5�g=*!�-��4z�c#�� )�Y
$�E*'�Re���al^+^��3K�5VbԿ�7�1mn�	�3��CBB�2������R��%پXo}zX���a������Ԙt���]ӞI�P`��A���.�ԛ�o��R?=co�ւX���-}hh�,XRB����[_�niiibn�'��}��E�C�������AXV���C�ǏXZRqq�ݼ��Ԫ􅀾:��Ć��TB6����qa6oX�?e]w8\[���Z��Ef"�%����È6z7��=� Q'��+J�̈��w��Ѣ�5����y����g���o�������mpz%iXޤhT C��1Eb>|-�)��yuǷ$�$���aٶ�;oL?f<�89�s�K~c��$=��8���ٵ�<{1L�R��|�bq����s �a;܀b�3��Vf�o�/��{,�O S���ᣉ��+�"��}70���8�sg?ȞD��`٠��������`mA��k�s�)cmk��ޅ���C�!�U6�}Cc�����5�5f��n�p�W�<Qk�(L���Ğ�拾�2��'���T���/�k�c����++����0ݲJ���N�0�����u�]�tA�����zF�}�����l�����a1��6
�"i;t�+[ �s�/kiiYz��v��JK'�$hJ{E��Hڀ[��3� Y�寽˾$�d?�Q���&���?�Ən�y�G9�W�{�Ah�p��3L�r���U���L�����[��@�G�jGw�<�@��Iº�V�[ fx(��6��+Sw����	��:��t�R��f�ӝ���s�b�C��!}�)׶�N���K���s�'�r�t�vk~ݍ��D�[��:ԣ���lj浾\�ND������[K�WZq�v�����$>g��}�<��(9�n��+��m|\�i�:�2�t�U�d�B��V��xe�J� Za�h��2��#�*��_��4-���B�5]���1�RٙE�0n�^�V.��o���Ŋ^]�B�ao�7��d�'I�����MW��	���19f9�]�H�^c�$ד�����Rj|c�����o?m�7z	����و��
������@9�h,{'=`�"L��Z�/U�z��u�G[۱ܻ��n��%m�yy�p��?������~��e�5!�MW��A"������޾dJ�z$m�cY�?Crbgk��݌�ŉ���k���	??+�X_�� �)�r��?�c��������&-jW�	CzBKB��"�a����@���`�;/��vr^q ��= "]��f�W"���DME��ѯ����7�o����u������$A[�4$��[K�%�K���d�䞈�V�2^�	&�Ϋz�����aO�3h��r��ٝ2��:dC^sx��6�ā�D�Y��4�A"M%�:�N��^40ֲ��#[�ܿ�+����Y�69t6w�X�V`=�ᰠ�UN��'g�u�;E�	_�E��~�@����?�����������>B�����8Lh�G&;mp�G�OM՛����V;�KrЏ�)s_7�}{���ￕB�7����P��1D�?���Wf�gr+Ɵ���~��(H��'����i��a\j���H���Oލr�Ƒ� WI�&(J�a׆�J�����mhʂ���+���T��I��&ݛ9�^G[|ڸ�����a�y�+�w�x��2m��	_��=FA�o�x�̓g��=g`-�Plr�?.��/_TC�U����kֹ>�c �37������*��V�y��v��Ïj�F���w_�8��)防O�GM������V��m�O{�Q��w�����B�,'�Re�A`:'�O���r�{��`,���w{�ϑ���(���;�M�"oi���FV�Q�$�/��3.�	p�1}Z�Z�lM�vX���è�^]Z}�tx�:�vr��R�~�Ǆm������|8~YYY಑tg�3���`�u��%k�f�s�~���ԬC�31i;9I��g?'���b��tM�5����C�����!4zER�_���T*������Mɼ���J__��{S?�6��D�Ӌh�k�*3��μ������#Y��Q��0����lD��iSl�#�o�:K^mzY��|����7+P�PK� ���������wi(���l�?ddU��R=7��cڈ/1r��+]V*��>Ƌs�7*���:H�-�S����KmgꍣΊe7���G2�J�
_��'��ѕ3�wߓۀ����HK}��իӾ�VA4u��B$��e�ϔ�K��>Vy@cA>K
��R��ۡ�{�I�T^p��d�րb�w�&�TA�\O\�BMy��LPF'�l��$]���S��f�Ew�$*
6+F�j;��Z�e6�����I�_i9�)��v#�*� exf�d����b���������ʎ��^B3T���[�v�y���Q�B��K��q>+}�W7�����?���+D{�7���u���[,���"4�.���#��H
��s1;3�m��IyI0X��h��E]7,lru��h`�L/L��p���p��7�4��؏��̊ղ�ߓK�e�,o`ԭ�eA��@�%&QE�9<�Ӳ����ص�ai��P�e_s�G�O�BG��n��X�ӄ�:���[�bX1.LK灓j5�qgVf�Jw��x���;
���?L#_e]@|��oـ5wc��j����%�+�N8Q�����:wR��v��S���	���TT{$:Sة̆����u~�}��8��u�w,��v���şw4��^i  �/��(j	��"H3����o^�>��t�������+�J�j���̹�XY�sXJi[�����o&�!�D��L~*3�c�.Yn�s���E�.�����}�LT���;�@_���wTz�����
�q��YO��7�9���#b([Ξ�9"6Y��8�/!���l�<�l�!M;M3v�	�����3�_����9ܾ�` ��ϻ��6�%��/X�9@�����^��LhjR�A"E%%i����M@?.v[LJf��54VT0III������S ��>�DOnn��2�-���W#�ĢMdV{|Hc��x����-`hQ�e���I��P�vz��e�%xlf<˘Y1��Nm]����^�ݚ*��)rs���h�Z���LL
���q2�@��vZ�g�"S4��:θ"-��0�'PdMbp΂�r6����	�Y,�meN���I�+SE�?a��ٮ���9	|$�y�yߪ��WB\�h̄ʫ=�9x-��X�F1��Ԋ��Z�vk��/��}�2Nh´�pv,��;�IV��<8_uX��r��_�Nl���:�^lb�������4��C������
���޳YT���B���a�[��Ү6P�˹��xs挠�r�i�vP^�}%�M0�fg��g_��+Rr�>CԤN�,�-�^�F��@���t�����ڔzC[F�Ȋf-/t���GQ��<����"�Y���j���m����ꨭ���^85VE<5>P3<L�y��4��o�ْ̧�M�4�������$��[ں�=����D]}�MG�m���'O�Η�ѫ)��� y�7��/z5tth��^�l<���D�՗�3*W�������8��`�6@��P!��"�ޙ���z�`H��H]ݚB;#(�{��,�n�h^�E�\�ʠ8�U|�Qc��%�*�����d�kZB�#|� ��<`��!x�
ryg$R�S�'�
á�I"��`](es��ς	�I��u7H���X�
�"t�*�`mi�����̯Y�δ��UH8TMM->))6%����zn~~bj*fr�ɗ�;�ǒ� �+'`@+4Ti(N�v��/o��[l9�����]zt}�:� ;X��j�/�–+�-Xn��T*� "b�e�ub>=L�U�jTK���C�&ߧX��q�&�IE+mŅ���m7:Vg2~��	��)��� )M�L�ᖀ�+����y3��0�����z�7���V�ma���/�5���7bz����y)b)�H��H�+08P�"]�~s!�;% ʀ|W��q�%E@s-�����?~s���ӟ4�=pc���O .�@޸р��L��T�h݈��1���3p����v�,f[�H:@�N+�s!��*�ס�x�d�
#�������T�Hy��
��e�y������RE �E��ʸ���o����o�E4��@�V]�Q�U��`����%���o�B/����r�ʠ)H�f��Z��6�Fd�`�1�t<�6���a�� PK   p�?X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   p�?X�'  '  /   images/cde853aa-4743-418c-93d3-ccba2bb5bc65.png'�؉PNG

   IHDR   d   -   X���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  &�IDATx��|xT׵�?��z�� 	I� �47�1v(	68�.�7�9��s��9/7��o���;n��8�����P�*�k�5�3��yk�33*����w��u����U���>Ҁ���'����eTT�,l���z����i�������um��	�V��
}[/,VT*n׬V+|}<���
M�]hj�1"����	�iD�ޖ6�h-�=�\�6eB?����#Z��٘_.4�z� 4�<M�h4���Lƞ2:ޠ������`a���K���ha:<ݭ`��4��S�'���U��l��Z����#<��^x��Ό&�Q��I 6zJ�F��	n$-vﻄ�}9x��{��	{
Kj�~���p�NZ�>q��%Z���b�현���>O<F��B[G��;���h��aC˽\�.'�>,$4Ӣ\[d$e]ʿ����+��������!:�AT�����t�J388��%K�����pE{���e/+���e������S'�aD)�7�]t�0�[��.w�X�Է���KO3lAh��O�ۢ��Ѽ�đC�
��X�L�b�|��&��i���c��.?���N�!�Yy���=�{X����u޷Ѳ/o��{�in�Y�n�me����m<7zf�um%X/�Um�3t`Aƽ{��[3�Ͱ��Z���`�6����w�`��LG�����E�F���׊�5�{�������~b��iAyy�x���s6a`�Fd!A�ĝ�@xR<�����8��k� 	�fSA�ރ��kkdL��55u@Mc]�+_G�ƴ��m�,I�T�#���T�o�w�b�V�c��U�o�0��ci�}ro��'��?��R�JׯrCG�A�W �q���Ѹ��i=�����|B��UU��������OO��x�嵰���|�0`�~��d:~����J��A�겏�,?�r%>��(���m�nn.��-��M�����N�߾�*(��$7���KB������(���n��f����U�G�)��94���}FLOJBuu�\���ѳ��F���	_�:z&��֮�RO���У'
���1kv
���c���#����z�4s��ܱc�9����<�b���{!�����,�Դtb��ӡ���'ڌ3��[�a|-Y��MCpP0��dY�V�����(**�G��w8w�E�%K�	O.6��5o�0c�?����
���b��igC ����b�Vqe������ښȊt��Qz~~>1�˗/G||����;s�Z[[�v�Z���)6K����e��'P�'eТ��ׯ_Gzz::��fM�9B��1=1��SH�������^B}c��WSS����ކ�!��4#���CU��h�_/5��������"��ъ/�SCEq8@��� .&��p����Zt>g�UV��	Q�Fy �n����}��@ ��S)�� ύ�ft�����#��2�����F�k,{x�2�5���A8��ϲ�hv�	��nf��7)B�(#8,b2w59�&B�wm?�j#jki�#���$f���0�c��(rk=49otvv�$m6���C�����~>��ҡ��E�5-n�Ї���� �܋S�c�S+�C��@b��� Y����4jn��埭f���	�ۼ6���z/[<ߛ'�v�J(�}���-���E�!���-�/%oЏ7�9��!��ȟ�Ͽ��H����?�!9�Q�ac_#�hd�b��� Ν��ꕙ~�=m�ԳX�IkGT��.�	��MKh���>�n�g��b���Ž�g�esP�`E�{��]�a��5B��<�8jΡ�fΞ=��������⅟�/��V�Ĳ�(���w���|̝3U׫�酻��QX��)����Y�}�b��i��XODGx� Y�ɬCj���u��H���}�o��o,��K Ƅ �`D�ya�]>hhQsCK�_�⃫�f+�
�j��LS�N�@�?04 �CΜ9-AgQf����u���(����s��Hl�7o�%�(--��1������@�J�/AkZ�)�8
��I���.��L���d��U4��`�IyMTԟ��]����sb�����A�_"����o闃�8a	T�PNC�5t͕����t\.k���z>.��y�s�Sŵ�Ƿ�{�ɝ�D�����Ǧ�[ŵ�ܬX����*��G�!1~
��.̜9�Hf���o��O�1C��ǊPXZ��j&R�r�}�.���4Q�$[n:�L��X�M��ݔ�r���H��j@wO�]�r�5��6�����X*k����Jy�AbM��.�6��>�QS�E�@����o���ny�^� � �7�H��F!��V��:�2fK�z�L�$��js
d���x�٧����0>���I(~�U<�%^{�+
���'6��9�j��I����%q����P*kZ�����X��w����C����ڋ�~�-}�����/��K�j)��c�"m�w��=����߿�Gbr+XOXӾή����H�p%�f���[��L�b�c"�-]��R�Ͷ�bE���bǩk�ĉ���[k�����f⅋��w�E�M��W�R�r��t�Y CC&����S��z��^A$V��޽Yҏ���n��=H0�.h��fpt�T���%����� �`'�����ƹB���i+���C>�0i�Q�}�y>Y�����(��C�:
�ވ���[(nE�qǖ'��S�4��@��wv�Ԭ&جF�?{{5S�[�sӹ�/��������	�1e�@��)C��7�k�����.�m�%�;:�U�^��R�W3�1P �;g6f$MGn�%�ڽHII&���ke�����cڴi�Ý�M��=��3䍈)Q�yy'<#�X@]��}���йhp��A��ة"$ψ�#-�g_|�K�ʳ�tM�+��M���b�CF܍��Tf�����E����B�!UWi1���;V{��:��R9�X��J�M��B��d�pZ�C��N��1Է�rýC#�2sz]����9� l�;��h���N�bˆ����������lģ�~�m� ť�Ĭ{���k��%��@жQQQ�q�e�&�fӆ�X�z��:"������ｅ#����/OI&<��+=O}���K \�(O?�����I�B�o��@��@�G��782�@;GU.n��6ː0SE�n�'���y��Z��<¨�s
I$i�����>�,�M��d�|�����b��0okx�hn�v%MHHP�[
APp(����5�ITA����U�Ȫ|s0Yrep�����ic���۪�?������2Y4��o-�!���,�*j�ʠ�d�[HH ڴ� �'�ΟD�%�� �\��˿�wDDƐK$a�5��e�����b�JA2�l�A;SY^�P�|��\����߀b1*z~��Tb]*� �eq�SewK*�r=�`4[a m��V�������v���]Ӽ��kHJJ�+0TC��on������]5����I�s���)G�3�d�9�,�3���q��y��S68d%�r|i�>w�KýK����=��%4ޤ<TG��&�#V�պ���h444`�\���'��<%Oc��
��c Y�J�nR�K�.��\�ncA��ֳ0���d�����i6��!(\ppax�c���&6�3`8/Y�z�Z�������F�v�W�8�c3��b{�da���
���%8�sE�Z�}�*���
�z�nJ(})�4-8� ��Ôq�	J�^�V䴐��6��W�"ƙqhX$f.��(v���3�O����
��H��2�q�d-\�N�P�݅�"
[[��9D�?A�lvAi$����8]�(���	�oh��n��M�Z).�bǯ�+�)������GPP�h���7���8}��\�׷��������oi�=������Fs�D{k�����OBwAeu���A�4�~h=�O���:�7w��X�|>��E�F�����?�qR������p,� YF~�?7K����_�����>����s����w'.���Ծ4��ux��A���|��{b�bAؿ�,*{ wQ\��U��X���aгx�i��zK�(�Ήk�W5cO�b׍8wp��YX_��A���&�"�oR&��P3��ʕb��х�%����!�T��WA5���W��~�J��>��>�y������3�H?.0n��#���� 	LC�~g�y��!���"<M	���}��K|���YgW?N�u��z�$�!!���{`�J�I��T�j���LAY.
��xC	���#��/1GQg�X5�f3*��6��>h��zΦ����N���Ή�+���Lh�����-䭷��)5�,����������$wlhhōF1�s���
7k;�!��0m
��$��F�Gp�|||�:Z^^.4���Ӣa��E�Em?(O�EMn��.9�ze��{��'�g�b	An��c�F\���5J��8"�@�U� �\�3v���R��=v��4>",v��uY���C+2iɓ90��e�������5,.�q���3��"���Px�03~�Ĝ��F�x����=;�5?�LY�g8隔�	^���瀌�=)�N�-��sJ�_�h!���/�Ё�ؾ��-�G�ܙhl�CuM�,JCowN�.�$�qS}�b~�ɮ�V�9�Jb�Z��b�$��3�/�������pP��|� o_>�3\"�4;Q�>$�d��X@l�BSc-����ҷ�)x� ui��K�G��K�R�T�d*8�k6o������D~)
Kj���� -.���q��?JKq�r���-O��u��qqY�fDᅟ>Eq�{���K/����,���8&|��A��B�ł2c.�Yne��v��P�8w�,����o���q�c�����T�[��]�9�;�;	�ċ.��Q�Wä́�J���W�o%{�0P }���`Q�jY%<�*Q�X���=���� ��A֢ę�������/�� ��=��p�5���4i�ܮ�7�����[�p�,��W_%�Svv�q���C�f�v� �t��N-�[�x�u�i�#�w��蘷�X���2�L.0	�Ӎ�H�? f�=�������J�.����a\��(nG���+���� �Ƨ���Im�����:sN�1�:s�"�!��HI�����1h������q�N�Թ)����M߉��H\���-9�ėdb��� &b�Z�
:r�=&0�K�1�M���>2zn�ǎy�kߕ3�Ltaw##.�<��3xl�ZIƸ�544$n�vm�d���!�w�А�ո��y��!�qMJ��� ��ޅҫ�DS�����1�hi�Lln�}�~T�����߈���VQ/1$<���b��Z�R�t-v78s's���x�Br{g�C�k���G�H&�B&� ���NcO'ȍ��a�SP����8�dffJ^�?0H�0
,�ñ�HH�G�|\���ET�<�m�w������L�HY���^�cŊ��{�E���K/�q;Y�s���ٗ�������n� 3nC*�{P~�A�]�#�X�
���Q$����cI)�8a��j��RM���wp�"�!�z����]����r���kp^��f����%�����RF�Ml%��#9y&YN?ZZZ����
�,Ė�N'��x0q]���l9ƶ�Z+������Ϙ�˗������,^8Q�S���{&�V���R�e���ק�8�Z_%.r�'����R�A]�i.�A)�8,DkO�6�8�HO���m������">���Y|{�$�!/$���	���XX�mڄ��p�*�^>-4H���Z�W6�kye;|�#���VW�Efx���Cs�$!u">6Lvj�m�^���-���&dȒ,0^ ��S�̳[���qY%\�t)������,z㾅!���"(��rqQ����/��a�T{��(�Z����r�?T����2ZNq�>�[sh>oV�{���-��[���u)[1�S7��5l��������W˒G��C�CH��;�lQR�WY9s?��1lڸ����;X�r%!��عo��_2&-��\�����������g��p�}8G�ȍ���O��6�U�6�?��0c�=���s�u�Q���W�Y��h����k��$���X�9���V��e�G�n�7D �3$�u]��|�wE�1b"�I��cB�@<hMJJR���*��T�E���^���m��� �'�G�Ɍ��V���l�l��߲e�D�u7����S֥y]{b��ƍj�iq�~?��I��_|IJ9&%�V�����(��Q��+���(�ځS���:'o��D��	B���D��Rb�U����h�7VE(�X�y���8�4V>�=1��^��p���C���k��[ٕ���}��C��|`�<�bf(׿��:)�Tc�ԩ����%A��/n�?1����e�y*�;F(Q\D��s��P���;ضm�Tx9���{�xc^n^>��N�ĵ]=��k2���KIX�|F�.�0PJ!j%��iK�5��ɝ5�&B^�8�XY�陓f&F'y���[���(�1D��S��JA�hjv�-,:�J
�##F<�C�B���OC�_���]Ɯ9s$�O| �h40-&�^z�=f�d���.�V�ܶm[��E �S��s�l³Oo�߿ډ+W�	�
���B��T,��tQ����=v��~���6��ټ��L^k�n�pը�t��\FK��!�b�k׮A��w���sx������x����ąbF=X7twŠ��S4���|Ll���PPP P���H�hf�#�o�v�K�{�hb�6n�(��1O�:%ۂ6oތO>�/^Į=p�RYE���QqwS��G'>\IE?c�k��ǕA�����¢#D��v��&Bg(�;*5��$���&h����&ɜ7�>���j"ƾAsÕ��p��!�����({�fr)�?���Ʋ�b�Ú���J((���2��x|�ܕ����	����@j�0f!�x|�T
X���X��>J:c�]%�ra}NC��D�_�P{�y���fK���J��t�111�ù�D�z��j�Ze�O�cjT����s>�ck[8�J	Ǌ��h�h�)�H&a�	4�,��p_�uܼyS��k�����?�1wӃ}n����p��9����K�a8+ ���&�/�t�����;`� ����/>�^���hқQߤ��xx��wv�fn�\��1I���Q�R�ıYm��c�pcE��kW6�o�&@(����ш��?��(3w��ۈ�n�}�"0�ż
���?�C|BupCY��Qy������K�����Z=	G���:e��^��uyFY��1�����TRBy��
�̓�"���=��Y)F�����k��h�@��Ga�A�c�ю�.E���QRV+��M���x9^�X�r���p�r-!�v<�&����5�����I��N����h��Ƈx��
�O�$�<�+��^{���x��XY[�y���ݱbq4����
q�>X:?� ��,����.]Eiy�n���42
rD \��+%i�����<`1�R|���Nӏ_�x+.�;ػ��ɿ��$�.����݅߿�^��s����cG)L]��g�pa�HP�z����M��c��� �m�ŧ���c�����'ObժUξa�~�=��D�ux]�4܋�2�b��!����",؋r��F��|��Dc� b��,>�σ�͂�H?�X_whMFG��H^���h�+��ᮓk"�}�p�q�ǌ��1�*��}��g��Վݱy�6Vf�{��exhe&4�����a�e��3Y�[�U8s>�*;e�����hn�Ǝ]gP\xQv�\�V�w�y�\�;����Z�AB���p�y077WٰlG�����l/�8���������%u2v�I	X�j9�otK���W������u��<�X07��x����E�� ;� op�1S��u�F=ŋ��N���v|�" q��Xɉ0����q�7gf0	��\����SBQ^�%c(p<'�rT=n/������e�0����O|�mْ��7޼��|��h����?�I�v��R~��*���"e�Vd������F(��j���D���C9��o�8��{"�rrrD ,.rrܺz�*v�9�����7�\(9,-����.I�JJK����!�h�0�����@;Yi[�e7�p�h'a��u��j���Bp[Y:�-7�<z�z`3�p�J�@�~r��a���O�yݽ��lŹ�~�~3:��0@遼�g�V{�tn�R�xa�U�d+nTT4<t�۾�f������"�,5��a������o���`��T�~��5t͚5t~ ���RV�Y�f��SS�L��l�1�w2��U���N)drѲ���`�I�:�7�".�[cs'R�b��N�S3������ȩC().����k)���C/Z��x����&ÅN���ǿDĔp���_}���T�$@R���䋅�\��5�>wݬo��M������5_�E���ܭ�w�8,
�h̷�ٳPUY%[j��f���MG��e�t8]u�����F�f?�OA9�Q+��)֠���'{g�!8��!��M��!+�l1S�ɔ;h2*yÈ᫯�ܴ�+a��p)����Ņ眻y���������J�M�Gn�[��nNMH)1>��&"�ew��P�#�Q���D3��L�?0��(z&�0;?�!� <��
I���(B���M-�&M�hh�Ĭ�L��š����^^�a圛���gNIki�����'��#����XݻBG1�wG4��W�U鷼�梼�6lւ�� ��y0U�>gڮ�@���^9/R-��O�������<M��4���n��d�]�*���y����F��'I��G�j�o?r*����K�#Z���k�볏�s���M����N��oŒ6�3�x���Y1��OX�Ɏ���	���Y޻������*<;�(�~b����w].�Z�����\b��(��z�ǟ��ٟ�|?����ɰ�#��x�f�׮|rWɕ��Y��G�i�3o7�mCցKa\�[�&������E�76|�u4̕��c��Μ�l�墚;�.�UWU��֔Y1����=�r��m��1�{�] W5�z�<�s�+啶��Wڌ�W�r
E��-3#��ֶ�m�3�[��(�1Ԍ�Ľ���m2�,GO	m���{[���2R�-���6/m��[8�%�T�HH�(��&Xf_����)�o�����(�w��*���V�{�3��ڴ9��G�~|mk׶to����-#���ⵇi$ =�6���	x��0��2,�'%�K��YSmY��o�Hퟥ�#�F�m�')����7ζ��Eτ�aBcE�{y<��7/-'ϕm��;4��Et����ϰ�����Ϟ=3�\�o-L���n���`�����8q���W�s*��KM���ג`�y��u,����D��~��1�F�~k��[8���l���f8.�NN�w��m��0�����Wh��k�g̍�w�y��+��5��N�ҏ,(�h�����֜n��c����DS�;�mvZ~a��V��c�үRh���{F��l%L8�`��JN�;���/�/9PF���3���=�b�v��:��Z���S!'ϔ���·٬Ԧ���?M�8h��:�$�J��h_����>%��I�9h#i-��_�cp��Wc�-����9歚�^�� �q4'��j    IEND�B`�PK   p�?X$[��>  dy  /   images/d3938c88-0382-4189-a86f-3cd234ee676b.png�XS�/DEG�3��F��"A"�iR�Ch!JPG�hPz@E@B�5DA�I/��ZzhI����y���~�����s���yx �w�w�k�k��Z���i���ñ ���+� �}����J}�n�k��o:� W����烞��} �z������@�j�k�p�E���A�Pg�=\}��z�?��vL�k�@~��\�t�?ya$�E2*��dر:�e��T����wkn���@��Y�G�ö�7͋�'����+��Se�o�9s��T�Z�EFl��G0B�n��q?i��~�m�}{,�Z�ô�J�j���Vf��ʌ�Ǯ�8��|��_߯��?�ҋ������`Sl���-Z��{[U���Oe
.��O��|��5�׉�V��Rr���u�g8b;S�p���a���1rͱR��E2��ď��&(�|�ӡ�.�HQ��:�|�_ߨ���*�7?�qk_*��ʸ��~��r�6�1G��q��qt�:Z�����@y�܏�)��sA�{�G=�x6�e6�`y��y��>�)Wbj�}bZ��~�=;;c�*��X>��@�M��_��#2L�K�W"1&k��c}�DXd�g���yJ���}��U�;����)���7�腳�$�/�Ē�5��`�jn��6�x��0q:���7�#��裦��c���ޯ����y�\�4�q0�x���65�C��Cg�Ő�V(S��!UsJ��!W���qp" i�����j�K�,��9�ρ�MH�|��&��	�`�p���V���O�����ga��[���u������Do�#���x�-O�QVX�bK�U�L�L�9{�5O?,��~uV��]�%�������?h\)�Ȗ�k0�`�H>/��+r��=�*2����{���>�
.��ZX��$/Tn�S��3���|{y�p��������B�{E9������b��6oe�m;�J�C6K�7J�����J�X����{��E�9+���zb���&ƶ�{rڭzSN��&d����S7��c�r�԰���(��)�;���ܧ�'���W�v�
�3�tڐX.�V��E��H���S�y���A�����o�����j��>���R
���U���������Jv�S'[��tB�\r5�io�ȵݲَ�	��-�ha�̐٘A���$v򱎟�&J-$W�6������2M��[�:����\!��(�jhp\7wi�ȭ弹���\J;��@pl���	:Ӝ/��%t��**n��/���<���)��ؐM�y,��#g�Bóz��w��
iB��j����j��:�Г�t$����������p��+�rs���6�j��Ba��l�Sݛ_c6��t>"m�a&0k�\*�Q"�pML��+�bv|�>MU>��B�r9�CG���/z���儐�̽�|��;�:e��5A	�d�N�olC7��bO�?����>b���МQΉsCoK>�,�٫o�ٯ��^����TOG��X���w��O��L)�:t�"�Uq�k{��F��w۪�>0�%Ii���Y+d{<��3S%q~�=�Xl�<�!%��0[K6u �ʯ�;�f�o���ϕ��X���ZE�����\��m8�4�бy��d�
&DQ���F�k5��j?�
d_��#F��l�r?)�Z��=�ya�Q�պ����=�^�xY~�.���N(U��P��p�}0XJu��/�s�wX�QNz�I*�M �
*x��Y��6y$a2P'%ebI�C�(?�ADǣ�� ��eS5䗖��7;���&�?����_Oh/���}(��n��c��:Ir8.��J^�@�m+6�(2{x}�����6i�S�j�sZ���!�6"k�m��ǌ-ϣ8��B!���}]��3s�s�@*�o��4BdM�hx��n��T����)jm}��Y�R������@H7p�X*����l�:�}���w
Ka��+d����,�|`q�t<{��6ܲ�^H��\�����5�,�R���`ڔ�_��u2㈺�{Q�ʱ97]s���o^Ek4�Y2�Z(9eY�!tf�НW9S�p��$���@�ܙ�`���T��l^�w��(Uq��ʥ�ʞrF�# GE���p͝2w�t�������o0��#�,�@Xp��sU+�
"s6�au\_����I�~�5�<Wǟ��8�X���Z���3���,��X��EA�s������k�\�Ќe!ێ��M-��~I�M�(�<��IǊ�UW�嶈�y�j��O��lз�;�6���*�?��� �L�a����ڰ?v��및7������f��:[�gW�X�2	�����θ���Y]��xkRS�����܏@ y�4��cb��ℤ6�h|���6��R�-����a��hǎ?�+�=j��Mַޞo5nz"`Ϲ�*�Hjm�#*�B.M��k��q�uEǃtE��F��Qr�WTƷ p����!����g�Y����{>�y!�7����u���3�P�!U�*� )Vj�t�U��S����[��Cm�]�L�'�_
ǂ��p�h �B�S���T-5�XJ��X|�+�x�`���o���Em�u�w��R;I/�;��kGae�~�/;(l�u�"��ʾ?��Zڷ5�6�b���)Ջg4�ƔDZ��Ԙ:���Mh~{G/.p�����"�WNݩ/��^�M�R��[l����o�1Q�oU�ݩ8��GV(�rƬ�WG�d��MS�t�`�Ԉ{7���vTQ9��]�H�U��s37O�����Va>���K/����BN����Q�!�� ���#�|az-��?�SX]�r/4�Qֲ�����#M룣���L��}��h�[!/?���<�<�T/,��.�hOe�}�ꓒ�Y�p�xXy�3,�7er��!KL���c����#T�̝=�O<�"e!	��(���{ep�_3ј���"4cOJ�V�$J1��!nğXحe����Ap�&�Hh�I��#Y�ԯ7OVN�em~aJ|��Le%ҽ1/�!O��'�NF�	�L�&���&;1h"A��7u�i[�W5��X�<�B��
�\���	��.�p�\�p{���%?���x���xuS5�ɏs��ӹ4܄����+E�)>�"'E�͙!���w&�A�=C���;�f�j�,Nr��h߾F��{�h�D!��8U���A�۠q�w7+��]	����^k�&��\�KG��,�h�� ���1;2.�,�{���s�N�/���@9u,�;F�(x{��Y��Z���;9b��wkG�J9KV F������9k1�����;�5�b�v��էsY���'q��Po���ހH���|��_\�Z�	�[��4U�9NՇҀ�['V��E�D�W�F���z�:&QS��0�cA���,܎�~��Ԧ��!
��� �f߹ia][�����A�M2V���KTA���}��p��h��+����0#|f���x��v�	�KL�"�_��Q�s+�VRl[R$0�wJ�N�f���f7VQ��d6�;��ݐPI: ʍB�uscW�"�	����<^��2H �@��Zx��X(�7��[���X�A���Q�Ԙ��C<�p�� C��5�"T��-1w��Pm
���{o��Or%D������|]N��#��ꍴ3��X�������r������v���8��x�"p�u�m��B���Ҷ8�rm��C�����r�4���}�IGsH��Z�v��y_!���cs���#6>3�ժA�&l��u>-�6���^�(�}�י�KtJ�\I�A�;I���j%`�P����';.8�6G�m�<DN���6�l�Z�pYʍ����c�����b>~_�k�/|��I��1��E�;H\��y2zA2yqd?^���:[��J����ſ�I��.=��I=�~-�\��A��ҵl3��b�r��~�v��D��x�+�5Ǆ�^�3�����;ue�@e+.��N"J��#͹���t�
pS��˞����t�~�d���Z{���~ِ��e����n��=z���}2�aE)��-`�LsZ̅�̷��1O���m�hn�k��;��ivA��;�̴���`R�Rɀ�M��9�����,���[�+���1���2B.r=���?�����$��G!]����a�/�8Zi���[���1r�c�c�xm ��8H�ԽrR>��;s�׮�Ԓ5P9�(H��ߜW���^I�����B�⌯Q�h�5#Wg����J|�����5	�<�~����
�R/�����	�	��^��m��v� N`H&�?�W����=�~���`ҵ׮��8Q>����)J����X^|u,�	����u~y{9/�	���{����,Ч�3����=4�=ي^��_��� �r���3����o�uw���l��C�5�����U��|MP��ݿ#?@�n��O�����]�Ë������-=��5@qq�O\]�-��<��u$ew{���Q�)�V�$�ڲ^~�?�Z�"!���)�����v�."l�z=�e�R;NM%h�1�3��U�b~j��|�q�� �E�@��ȅ���BjX��A�t�]��?0��E	� �b7T�:�dWk�-:���~����/7ȴ]1{�% �$�ɦeS�8��k(v��v���H?[E�@$&��H��t�>1�v��(H�HG�]�����c���wB^��j�-�TvV�%�*XY�]��6��@mv��M��0��S*H_ݰ	���@�fo�)cY�0ⴌׄ}>�2��-a�N�Q�.S��z�	GL�R�*�sJ������<|Sh���6+M�T;��T�_ۋP�Ί�u�1����ɟ�jK~Y���^��G��>ܖ,nD&�!�_��2Z���TO��ȼL�:�-� f��]4Q�FX����������TK���ӭ��?gnЖb�^ŷd�����j�����kwrc�S�~�I	�ZL��dK<:83G�*m:�e_Ğ�`L/�m0��5j��Y�� N�
�CC��Knn�,��(�aϑ������Z��f���]��BG��5\��;z�܇<���y�z�j^����ʉ�Y|�Hu��i化��L�"u�	����>e�e����3�<����F9&��G��U����hBJo��)`�rE�>86Qb�{���ȨMMF������B}0���"���9���"�p���0�:q�BM�r�6�?~�y��ߡ�̌j�*���N���}���E��{��es���7���'8sivyp����o���{ta�:n��ю�5j �Ǣ�ɅM�Tf�D��iM�F'u\�#���Oܻ ��r�_������E�����/�����<���?��798�QO��;kZS��R����톻�"��3���<��>ʜ��ΖK�-����e
Z�%^���N��A����w�|si�=��t5]���l]<+�����ڧO(,��HĻ1Oa���G�c�/d�8����B���.�D����%�����X�_r��g�b3˥h��w��Y��۶5�ʧO�,[j=d��C���HyU�����i2a6+b�@���'��э�E��_JKw�*��BC��#����Ɔ���7E7�:�]����b�ym�!jXo{�ƟQ�i�R������چ�;Bܞ5WZ��w�*t�
=�P�z'p�bm��N��^aW�S��!3#�T[?�!�n�~^�Wݏl2���<�4�M�s��r ��<�/��=�)�>"�Q\эf�������76��GsX�A5�.Y�n��Gi÷��q����h1������m���)t��0���7j�L�|4uHɬ�p���<��\q�+.���[y��#	eϞ�æ3���~n+pN�>�N����J�S�4�[�w��Uʁ�K�aG+�Z�91��C{s�'�iמ�:i��A�Ʀ�������4��*�:����:KTԏS�����������K*9P��CX������G�Y?�m~�'��'Ծ �<r��;p�^��}�d#k!3�Z�ڝn��n�?k���A���>��@[�����"����5F���z)��޽(���_�}i6X�~�����(�m��`1xq�ۉ�3�A6�,���"eo��:9;!t����ם��Ǯ �pÅ����V ��rx�'q���ֺ��,J�X�)1x�k(�P^��h�B�c:q�C��u���A���p8If"e����P�%qJ�֕�໧��"���ɭ}�3t�4<�>�ac1�o�����_�|+��jp�%�z]��@�J45Qq�#@�>c`��r�Q4����.����$���yv�-�4�IUJ�.���Ѯ�8���:��(�ЇuWcky�g��I'��?ܴoLѐ�bA�p��f�6�m$�bxk�06�va�c�ħ�7:�UG8�v��)J]G�OY.t�vT�^��l\�G���a�������^ckq�����_��e���ǎ���Nx�%4���mn�ty$��.�f���Ӟt�mv����̠5l/3�w��O{��b�O�������{��F$�+�?,���˖��|r;�R�	����dO��&�Ǐ��zה�V��<�J�[(���ɼ�a�-��1�O4�9��&3��n��|Xm+���;������=�ia�i'e����ym[���qu�wV���@51W��u��GS����\>%�s_?Qq9o��BZ��Q<	e8+?�0����[���ﯱq
���-�%��c�{u�J��sF��Xt T��O=S0h�MĦ�4aWcc5Ә vw��������g1	��¬�*��mS�x!�����S��!�HVg~-^o�	�/������_8�|g�O��5 ֯^c����|u�c7 \a�e�5�%.)�����hvB�o���*c*|���l���o�reE�4$R��y�������ݾ��%�#�f�W56������`�M�y"D�Ž�'N���̊G|���P�������^ _93��S�dBh�¯�=Ӈ��
����W};��.�<�ix9�s��s�3�ࡏ펞;Qɯ�ِ��4Z2�G��~5�PEھ�Ҷ8�3����#��UZ~g�v�+�<�����YݒW9�`pn�b��l͔���\��M����$�<�`/�I!�T�dP���0T�gΊ�u�^��ʿ���/�Blݍ�������݈0#0O,8��l�~�
-�[T�[O�_�'Y�Б�r=���7�᩸�`>4	�����`�f�,�W���Ħu�3�0N&�Ȱ���?w��!�*���O�����.�*�`%�pUw���ڢL�Q+��?���*�H�y"ײ�n_O�r��??J���Q�|��a }�q�C8yk���k��A����$�8�[�]̩����Ѫ���Χp��ZfF�l�0>�Ϋ?��-��f}��o#��}���i��N�{$E$��C�AUh�M�Fe}��o��o#Vwz��U�{����&����\�w�sk��ёo���Z�R/xJr���w��ԟ�%z��m=�t\a�1���V���
���5�E������K#�f�/-�i~���!����+I�#��;�O��=�xEU_��������W��,�!�1�S�vP�J��t*�_�X_t��e��m�r��+L<�L�8�y�X�i�7�U=�.��ԫAӿ����Y�³f�ۮ�n^��Ɵ�ŝ����~K�?b�J+�Q.x�i_���1ZLM���m��U���K��@�굶^C8��:8���č����*K��SMǉ�K.�����*D.i��ˌV�y�q��\�*����n�C�t<�b��6��3'85���~,61WQ�ܕ6yR��P�C׀q�'�'�]�--�Ứ�b�j���?�U*��GA�'Ю%�����W�$;��ϳb�u4_s+���!�1^�Dst�ujr�V��݈��`�=���/��G)�:Bo�����Z`�q���zk%��2MK���u�0�\z�ǘ��u��% Ý�[S��|qB���|`{�P�mv4�V�G��g �[9���e�C�p�����P����=�3����@��,���$�3E�TݦZ?΋M�RC�-y��K��Ok.F5�����̗��?�OL���\H���}��~�55(#q���^_rJ� �U߬��uZ�cDM�c�5��t�.##���-�@jr	w��8E�g��9��؀2�_�G�+�O��ncrZi��
�5Vn�f��;Z�򋫯F�@��Fq2���mO��RY��C]���p����k���T-�H=�XR|�Sf��G��� ,c�68p�B����T~.P�cUr�Ԡ���ܟY|��W�V�Y�ӱ@��q�ʕ�l���z���\8���RnK�?k9�I:�.���W�C�+�����˄��W�,z#2����N��;��7��)[��__y���k��FA����b�������}�7R�O�8�>�Fa4=���zo�J�	�]�(���'�ޠ�M�pb���/�!	�����0؟R?�����j�!hhq��4��&�[brp�}Ɛ`�O� �0�L#�d5b�clS�P�V کYZ�\�6:��ȿJᲛZk���ډ,�*�+�.�gy��S
dw2o���Z�n����XA�eބ�K����Kƥ@���z��2��7�Y���
e~����>�����?�����o�0�"��!ic&���|IU�������:��o��2��=�H2
h�"Q�b���<�����d��S(8��0�s낽*{J{�q=K���џ5MF]�m�)&�(��AbU�TR���n��]7�j�����qI��
K�-���ۙ��ên	O����0�+:>7�KbF�SU�O������ȱ�uw���%#��[v*��/���DW��%�oWQT���/��Ш���LJ	�r�!0����H�X�ϯ)&���|��Kq��n�?��zȁ&H˳v����/�\��	D��_й$���S�u��Fͼ��7��H�u�t��s��2,���j�}��\��k�A`�./����V�:�
f��\�7���9��	��3����C�^w�������V�����xl&�c4��#�w��}8 g��{���sz9uI���zD����y6�cWR�C�GFff|�����4g���ޟ�	�#�>%a��o�TO����<ژ�n��9d��v�m,[�m�*v�H��3��1���e+���.���"�T��?K ֺ�����c�+P��"��H|���ȃu��KY��ML��8�L8�A�<�[�{w�S�l"b�g���J�I�z��O���M#���*��2znx��?�V�p�:4~*��� +o`e�h���~�81	�F�5=��,@\�ҺG3��'_%�'�'b(�@�)�J�Lx�����]�=����v�͒9�"�&�5��i�z�n{��1��v.r�V0�6`�x����o��c����[�v��c�O��C�c����\�6� �M��!9I��U��N�	�E�N�)Y�[�Τ�K7�4���K˛߅��%���C�Ș���b���+��Z`�lm���9 c���vt��kw+k.���98 ��eyIɤ���kYY`)�Ȫ�a7�����W;ڵkυJy?B�".eœT�1C�����E�����������^o ����WÍ��l�k��Y�Ͳ�_+'WR�O"�N2���Hp�[��an���G{��V�K��s�E6�M)<K�P��f�߰ tqC��=/D(�뻠w�n ��6�o��� ��*O����^T�Qsˊ��=���ھx��-��/�gA�rH�k�$y��}R\��UJ�~��|�' �ƪF-�Ƃ�AFѲ�nEՌ���?^z��t^��2+�V��s{E	��+�c�#L
l籬̔���e�?iK�N׸޵��ؠΦ��J��Θ�!��OV�؟tR8�`�E��'�q���%��Gɬ���:��S{��e/��'4�<�֢��"{䵉-g��V��,y2�sa��ׁ��M&�3\�g3S��Α�5�c��?�ۿ!�C��d��R9�n��u��G�d�gd��̭���/�fdf�P����U�4�$����C��/�8�Lp}���l&&&�%Jp���7�3�@�Q�I��N�$r:��n�.��{����	曶�#�7�q�fg�l/^"����/ m�Î�y�L'�B�D�/�[�cF�z;)��{Tii�.6�f�m���hÞv�-�h2�����
��Y"Q�����(���}�c�HO���$ ����X���Lr��PV�w���j��hH� ��,�#�r�Nk`�R�=-u��f�^ԯ_��A�xz7�N���q����k��پA��Lt��=�[����]9@W|�G��ىQMNҿ|�}x�| �5ie�v�r3�[M����"8v��^���~��p�6���y=9g�h�v���`j�]6���	"˓��u�d��_�G�͏۟���7U�0�n;���dY��wiȸ�+k ��y������=4.��1��x=ڽ�_w
�b�;�פ���C���m���e@l�w�*v>���I�~�� �N�ݿ�;�7�0.�}��<�֥��>����ޑ��$��6�����P�B���&���kC�3Aa��X!�b�$ʀ������M۽?�I���ϧ@��>�5$W�>��P&(�Ŵ�B���=�	�@B�-�U3���h�b[�4�)(u����;K���-#�I5/�,��(�C{+M﷞�	w���&�	^��wq�G]U��cj4M`׺�ߕ0�x�}A�j�\bŴ���<HH��6ݭ^�L�9��v��PZR��	[5@ EU�2���j]2gZ���`K3��Z�c��bK�.gY[��w����|�7�]�9�==��*ItD����t�5.Is�P���w���5Kfsx�ķ�]�$��?(u(��ȓ����^�z��@N|^UD[��4�C4�i�ɏbpר�S HV�x������a��	ɸ���c�)u��+.���?j��έ��>�x�ؾ0o��7vAC�D-��t�X�I�*�:}�[�U�H��g�o���f4,�����׏.�ӗ<�Q/KwEG@?��Z�t�SU�t2]�t�p��$�v�1U���~ɯ��i��Z�Ѡ�|f"8�
e�\c�)y}B����$0�Z���BQ�!��X�D3�Ȃ�G{]�X�LL0�Y�'���(X�tFG�1�[��l���2
'�%[6���I��7�������-:�M�g�c3`1=�n�:�54��:mޤ�`�y�Ǭ������E�:ߵa9Ucҟ��w���^p����=����N�X��\�/���N�H9�l�f8�c�0�]�����thdl{����RTWO,�]��A��~������"���i;P��t�k���kZ�,V��0��ʅs���z��YtoWaȫºޓ��˓�Ę�R�7�m�g9D�����{V!�%���0}�
�JuFf���� �7��m��J��L���ܰ�Z-�I��]̆�V�tf�������]���X��r����74��na��BnU��\5��;CTR�cc�p��� �n�3�� �G���?��~���Q�ι��ȖZ�w})����vBD��{���'2�5�&Q*��'�S�������M�*�Zr7����_�%�V�T����NVK�,^֏����Q���Ȯ��Ɉ8;�xZ*1�=�Б]K��4�n��Z	V�1��Rs�g��������O�=q�����d��dܟ5o�m�U�^ur�#U��Y�>�<�6�m��[��o_�޵td�� [y掴ʤ�f���$F���U�,�-�K	����ȟ�u���3G����>�����<�2�bu����sWf�r��r��t�f�`@o#dK���견j�Rq)���4�/�S�瑁v�eځ����fB����*�.�6V;�#��/��Փ���嗊�*�H�Fh����%�M7��=Z^S=��J�k�ȉ�K�r��hK�%O5�o��;*S�6u����Y�����y�*�������S�b�q�n���X���/�imRK�0La����մ$Y/��@5���.��Ex��)_ŋe�9�z�1֧ђ{w3$J�E\�0��cG4vO�������w�w��o	����s����@R�}�K�[]�Po~�)	�S�j�ݗ��m�I��21�#��?r��`r,���-�z�id���q�n;Ό�iJ��}�6��8�X���@w��=Y�`OY
Zw��y$���D)����?I��\�UP7�u�mIa���l*T{�s&��2��Wu������ȦKt�Yހfl�I�*p�b3�5vb���-^m�ؑ�̢����i��ȼ���.-�ZA�:d$%��9���T�ͫUA��"���Z/�5�I��;{��5�����Lz��G���4�Um���׍��O ӣ�
�
Sn4��g�q�N���R���7�K�(��,
�ڋD���ղe��⹶���_H'��fl��9rף@��mtT{��܏��˻`Ɵ9{y�/Q�ti���LhP83��_�
e�Ae!��p�����oXe��66��9(7�,8��A�Ճ�Б���Pj�{$�C�������~�NQbf�y����� X[���xwP�,�K.wa��l/`B��`q^�W�Km^�O!^�U�AV���lE��-t��cWq�rZ+�#k����V���Z�T�V�!M5!�����[\SzY�����[_h�?7r�%�ϯyۄ�n�0<��3lKSx�<�;��~����4�6���-�v�AVcZ-hc�)��cb#k�0#���1�ۄ(�I�kދK�I��/��]��C�q6cʞ_ͼw���R��(����=����LOR���M���F-A��M0F�ҟ��a�*���mbϟ�2�t�����;�E�2�8��p��|K��zq�&Y*%�?�ߴ5*�����֕���ï{�2�S���/�z���$cG��'���?:u��	O����ՊمK��u��8>L��h���:!��=��s�7�9;|�z쪺.�0������HV�����c/k;<H���T�����g	�� A;08���-O�?���>��{�0�u�	&�Tq���Nv������t=fmkXRU��۫*�
}o��3�`'���RY�C��қϏ��|�p�!n2vSп)�;flL�����[}�[,�YҴ���i~C`<�GȣVͧm�پ�����/�gjt3��NX`2硊��ͧ���v����5$o��sg�ԝ:H/�J�]N�m��8�����h9|��o�LWB���O�tn�h��:E�0�� ��Gg=o�n�ǖf�>~������ϲ�WՋ�֭�I̷x��@7�[�r�f�1K�rq�Y1;����5S��P�F-�y�e���۫s���$�o��`N#�������{n� X�c^DB1����C����g���}_kOs�����b�mT,sg�&^T�6 ƌ�*z:��ݪ�(�����������U���,�i�K}���.X_�of+O���cO�7'�h�{ĝy@͞O���Se7k�T�"�b25W�X(i:p��Vա��z���ɣ��I�}_����)V¤���e��ysp��0QAML���0T���o�wrK��~Z��i�`;�MO脸}�ች�V
}=)KE ��MيfwQ� qN�0���*X���9���]�d}"��9�>�H�\��Oc\}_�}�'v�-��b�&N�UL�E�R�G2��lb��<d	��J�����;��i8�9j�$k��Ѝ���B�?��$��2H15���#FG��k�P�<�y8W��T�i�l��0�b�i�93��4Yu�pϙ�Q~W�!S�9р�����7�3�]���$��P�9:�h��P��.r��8皻?�0�I��E��ocl��з�V
���1#�D�;~�P�൵c����K�.|�ϟK�/�iu�5��kk�'��9J^��	y;å;.g�d k���k���I�wT��'D��~�]U\�ՙ�(v��_�}�	�|�����XfS�Ǘ9q�1��D�Te/�;e~kb����������MA�J0:���t��2�1A�{���>G`��� -�D9�3w��>|1B/<�z�L��L ⓟS���7�a1�ɓM��
��֧��k����q&��?���:���Ji������s�,@||�p�s��������s�e��	ۚ[�����^�e��a�dW���қ�Gwz�����E���|���!��*��!�a�h��j���IN�v]P�gX��ml��&�u����hm�3U���h�6���@eWoy� �Z���7��Z����u���R�1�q���3��~�݂��������7"@$�Vc�(��A�礴&��!�m��B1�;7�}��>Y�P�f$2T"M���k�m;�vPȯ����Z%��󬱒ח�\��x���^%K�\?W�u��v��zD����
Ƽ'�	)aZ�C���w-ER6XR���Q_ �Y"t���GɅ��qӹ�;��0ݥ S0���5�P[N� *���a1�eF\� \���6;B��W_�Oa&P�m�XD�
��$xj�W׭E�;������N[��E�{���pǶ5�@�g3,Ӿ>�^;5�DGЬB��H�Z>A�x
������}�5�����U�X���~���=jfZ����:G�jX9��	�V����t�ң�] �l	�a�x*�,
^=a_-���@
S����i�n����H�]��l����!�BD�Vɓ'� ��U4np��f0�-��i*K�5Xv�	�h�</�o�c�x_�kLйfWò��J���U\�h�I��U������(*�a���TL�#~��B�b7�)Cz�_��h�2�����|>Ɛ-�}-�G�DYn�͟+B�y��'�p`�cp�F�_g�R��WtBN�8Vp�G���S���:�>:e�.Mx��-�M�E�ڲk�V���cm���շ��\�	�EA#ȑ_��O۸1�A���V>"��	/p0�X��J�K)ɯêc�3S\�ոb�iG��W���g�ϲ[��3���s�D�3��d��Ϟ�TC�RI	���Y{�]V�H����i�7+M�����-�a�J���{9/&�cJ�ԿL���>OTm��o��b}�WlV�D�f���C�����p\�ӓ Ŕ��m�JuoFJ=�����;ױ�ח�8h��:�	Qm�\/"����N�8��g�LH�����/�)@GIU���Tsq[wξz�v���P�!6k��,��]��W�_6@�9M�Cw9A
�(��ӓ�����ɵ������Z$�/�^�@5�EwU���B���=���>
�.NePm�*ǟɝE7��Km���C�c0C��n�8e�����}5�v����V���0)۵��4��pm����|�W�8S�����9uIJ�fc�+;�0��9P�N6�"v��x�U��rz�<�v�h�+�_%VQ�T��{x��d�0�5��/�_��U^}����g��~G}��D�*��q��;:*������LJ���wA��[����D~'|'|'��!�r���^���>JH'�����7]<u>ԩw���x���w�����d��τ��������f{�����k���3���;���3���;���#X�	@F1�&BR�L�xukk��&5! ��֏��ډZے��0gŌ�r�.ܝ�����~}���ESC���s��C�G��W�~�}�� PK   p�?XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   p�?X/0�m  `  /   images/f42dd85b-579e-4617-aa27-44ea24c5d2de.png�yeP@�&�H��w��]��!����}qw��NX܂K��x߫���u�T�t����twu=�LG�(I���������H��k�w�C�ϣB��w��$��
C�����P_$t��qSw�t�4u�����d�q�s�j�d���b�u!HC|.+!��}n�@���ftw��[�dk�}� �����J@LMA ��s	�s9p��%���Oz����P��&��``��)��<6����!9F���j��܋�Kߍ���n�Fqg�Y�j�Q�k����,	d<�� ��XX%��PB���&;�<� �C�B��}�D3�#<<(�&0�ߚ�Rq�2�H>7�x�?!���6�5��<x?j)�!�YP$T�Ҏ٩&#͂N!��lS���T�^)Nt�헳e�p@�^��[�S[`��������|e�#�A�gY�n���<��h��N��.��)�ʝ��.���A�lw/�\ʗ|بp��V���1�ߞ9���ТJ?)Z"8���<���&�@��J����P!���w/�60�լ!fI�v��+p;���mn��=���Q����z��i:���b/LB�ӓ1CP�UT�
(���b��(Ɇ��������T6Jp��=]�����$�N�u�A�dX����]7̵�R�:��c�;iV�@�!��B������x����k����(B�c�,I����?{���׉�7�C;`�C�O3��/��G�/K\�X�B�Fc3�	�f1�A�aj5b�dL�a�嘢qxď����'<W��b,I&>��SעK�0�N��e|�6�_ �gm���~;;;Vo��S��G�^�ߔ�G�=}�U��љ��J��hT�1C�{�0���C�&fa&2^�A�" g�/��C[l�p
Y���R�F��lR�.��,�� �	Na">?�7�q��Ճ'3�u�O�r�/��^f=9�,�F�s�^ǧ5���h����s�_W����@~�n{�q�\Ȅ!�'RS��4+mk��ͷ��^��zx~+F0��
�C�F����E|rz!�l8fE��Ja���~"�����q)t�Ŵ��O8%�Ŧ�2�b��>��8E2���[7GG{¢(A4ɪe��P˪�-#@ �	�A���:D�T72�x�>�d��&Y��2}`c�!����lXa��Y����e��� &i�	:�J��{h��;CO}�~+F�7�����yr4������WG!�3�_�D���+F9rѯ���βh|E���4�ޟ������v���#����g~%���n��Գ�j�����W���s��pa�֥<L�Im#>Ĳ����)�@��5u
��������{A9W�M�DmnO��<���5��Ā	_�o�zt5s�E�F�s+�wx���c~�]��ǐpJ�{/yڡ�Þ��R�?SՆ���Z6���I�B���R�LF"�Mbt��)y1��F�1=B�(�R����/=���T9gU�R���^1�mR|}�Ƣ�/'05�Ie&�;l��)�k��/lP(��^�Nq��Ca	���c�g�Y{�PSS�t���#ok��T@��H턴X2�b��66���bKGvW�)%@rJ��--�׿^��[rl�	�VcLU��%����.���m^��{���C+8UH��_XA���Q���9q!I�����;z��߃����]��aa%崛!Uz����ˍN`-��S͚�*����l��M� F�-dė0�&�Ljd�I8�!�L�C2b�Ȯ�޽}E��/�}�?���'�Q;��k��k���;��Ms�4#ꓔie'�s����/e���ȸ%�o���}Z-A��KcO'��)ö�����fT|��������<+���N��9_���/��3g�(�qX���5�5��!E��]l���g�[^򀉪/!p�Ȱ{��,�CY
�=�[Y2U>R���i:&@C����[�*v�+'����T��t��MҜ���H�����`�W��Oe�de1�w�m�З��Vf:��g������:�5!v�,vX�"�[�)�:h-��k*��+X>����o���x�h'c�/,Ϣ����E��?j�C�e�1��򯖹8I�|X*���6�	yD��R#��%��7f��y/ø~�K�2�;��g�R}>*��i�S�Q�sHƳ�d��.��h7@��֤�Xw���bFQ�����$\�GQ۴��P��d���Ϩ�'�7�Z�����msZ���O�~��{x�ܙ��Tw�ոS��c�(hNn�N�-��6�(2:cf��qmpQ��>]�Q�М�]��(jZ]�"0���$�"CI���&���Wt�W{��"���7]ڳ�&'�(��
�6��KU�4E���g����f�W�.6.�:���d��,_\�,�X^��A�\�_��PZ��,��j���A�~Ejk͎��q�`��C,^1��w�F�?���w˺�Z�����u �h�~q��ZͲä�<ʮO_���c�R,�+�+��ٳ4�Ֆo�T���.���z���(@�GU^_���
�1E�����;����W�nr�N�G����	���X��	2@	1��f�I*�?�;�a�q�ܘ�����,�!5���C�d�_ڮ��x�~7$�=�ήf\�����&�l!D.+E�I�k����z�\*���x��S�1�i>����T�W��!8�g�ɻ�4e,>g�=����_S�d+�i9�w�a'�?�%��q���k��2��0��YK
v~V��Ll���Tx�L���iKx�&�q�R�#�_A�ߺ͊J*�ݼ0��/�����43�����1��t���<�b���K��
n��\:������x�\�B(��z�$��F{�l ÂgR��7Gޯ[�R0R�u�l��T���J'���r ��3l0.�b��}]�3Ѻ�8Ls��jAvl���g��s�qH������9�{�.��4ި��!�V⃪ߞ��嗓��¦��8�`�h�1x��8��'8DM9z�]��$MI!!�5v��&�I�2���]j
��O�FFEd���$R�Oद�ټ/�Mw$��X�u����ڬd2��b��Dՠp�TK��;&��Ω�~rl�#R��WS	��^i��]��A���;|a�퀽�<B�_,��_d~��u�v�03��A9��Y zY;^��Ob�� ��=x���Nr �yI�b��mG+����\�;��=2:<j8�[~8�]n$����T�����!:v�	{?@�;hG[fj�ͻ������o�YJ8�p���|�i�=L����|)Uq#Z�z� I���T�`�K.��x�5��y��5�s0`��HJ^ȉ�)���ݲ_<S	.ӵ�"���;������1�&O�R�5� {k�g�sr1��;	�tE\/�LsK+X�� ��i��U��;�.��0L$U��p#�GfQs��,���U�����y;Z�t�>V���	3��x� ��|�Z���RM:Y��|t�h��>�F�$u�S#s\|`��9���y#A����^�W��$]�`�o�"�(>}j�+�bԾL��ו6^e��5n��̷����ѐ����_E��l�J�}ؚ#o��R��uv�;'�{;]�.���y�P�L薤n�-�axS���)���&� ����;��CP���	G]}�ձ��;�]6J��7;�8r���π��q��O���ٞ=Z08}�z��I9�����a��+�����-.)Za��s)�͍�q�稧2���;t�I$���b����.\BW#4Њ�m�6����]Gg������{�=��7�H"�M3c*]���H���I�R���"�T��j:�!�yga^2����)ñ�C	�#	��x#z����^�G��[/>��F�����l`�Ы���/uLE�f��X��;�����)�QY~��?~�k�l�m�I��$j@-�ڐz� T+��31Z��Aaݗ1r�����-$^n��G_F��md2ø(t�r��-R���&��wl��I*=2���N}]��Y��~�N'b��oɕB�'b���ʖo��'4A�'�[��ވ��w�Sj�FxsC\f;=�[cNA	"=W�@z>;7���� �vѺk��W����w��0��B����@�u\�hٜ��3���Z���p���%���V��G(���h"��Ȏ�1���X�l�����g�쾠��:��T����=AWܐ�=��x�C$�Қ �&�%�͠�<�Q�e��n* �o_���{�����>z�p��0��w���6��81B�v����ʮ�/��o��;͇�n±i|�/�6����סiL�伋κ!H������g��(�9[7�6R�*�D1ku�Iw��l:�Ĳ�5��iJ{8�s��Y�a�WF�	�C�8�dGc�.��A\�ߞQ�~7��l�t�Z~Ϲ*6־��&������\�j�~
�cpC�U�og�uW^ƻ�Fr��	dK�D��,�f�%�`��[b+S�k�E�ۥ26��,=\k��P� �l�����A�V�s(9��\�p�v�=���/�ֻt�d��H�wVDw�+���j��Y(�M��~��+����cv��͙�)�z7l:�ӛ#PL�B����l�0���pE	���&#�����k�< h�{/��Pc*�x����p�/�����;"+�)�.��u�!��hQ���c�A����ȽdS�A���'��|�+�}�@`�i��! ��|�6�^���#�G��[��AI�L�L�������b��Z6fa�d�_�=k�9�q�s&fp%њ<~��9.������Dr�b*�O�) ���	�*LH�p�-�s��,͓y,`��ж�sR���"	L�R<�Z�Rɡ��	�*:d �T���P�d>�� �=$��kwGږE�upz7TM7��޸J�� �2>�@�	��� AgX:4�m7�<P�t�i}P��5�$��
��LMtY�я�7'�	)#}��{4�f �3�������A�9l�����MR��?'��Z�s�Wf�FǺ9����Ld�j��\��ƪ�Tc��f-uW`�ѡ���e9��t�ƓS�aK�
�}�.�7�a���}*U��jy������S�#9�S�>�DEҟc� A_�o'�gm�������dR��c���_��V���O�`,�]K��%��_~8n�6���H�4�M)�� �?n��U����:�j{�<��GQ滉���koP���v+j��#[>�����!�t�n±�+̺<�ታdKGJ�]4���nG=��D��{���
�k<�z�����Z�S'{3��?s.������XE�9���:%�}ڃLd��KUw�����4���[�:����]ŗ.�jq����/.����[!�,z��Q�߱��B�Gr�Z�*B����`�ۘ�|=�}�Q`.�$�&��Z�v��䢕��!{,;Z�A�ȯꠕ�O����3q��;	j�R��\�W�n��*g�'#_ �8�a���h��l�V,|&_I���#�;�D�<�4W���u�=T�|��λ���|#��u�3��t���"�8e��Yq`x�h�}V���.���zA�>��ŗ��8�y~]�8�p���S�I���ߏ�#�S��.����W��1���N�����%�0����=V@=�:L0��ZGl�Ⱦ()���`YS諯�U3�)���2ʠYt�#{ۂ7�`��?h�Mn�gioi���(�#�дJb��f�˓�ln~��ƫ��&~�xi(�o��<~���>TK�L��c&��œ��aG�k��TR1�s�j����B�ƽ�^R%�x�_CK/�r�}�?����oQi��Bf7���(��U5��i�L�R����k�����_����X�W�Y��b� KFS��$�U��<�-ƒ��X�_�BJ�o��;m  �B&�gM��r[�9�f{��T\3�i�99^�:�sL��j�qi?N/B���
�c��'�D5����xG�x�zt )��֑�^�p�;�ݧIS5[�o0ǵ@�x��m"��H5��[Р�gN~dw@Ҏ/N��lu�9F�*�^�GF������]��P��0Яa{��u�;ɫ�5��/���4��m	'/5g!���V:���[�����������)<4�K����ƯXSn���B�����*�4|�+l��E�2�9ڵ�����i ��#�j�dD1�YIz-{�7so��:��'�����p��`d^7�#}���"�e����ci��ｵ����l�ק֣�
<;ϻ������o������1[��.8�4��->�!I�ܙ;>DHY֋%�:8wM��@WtRR��?�?�nW�}on&�ȍ1�桭�q����/ۍқ�������nLeO	��>�ݼ���W�)ӧ���� �/	���F�eG�F3�%V������i�]i��]�y�n�A��0�^"����_��װ�3W{j�4;�#��	� �4w�[k�$~	��'�1S�M���xu9�X�M¡�5ZEr-C�g�c7���u���z�hn�0��~��K?�wcL�P����hv��b������n�N�&{��H����ӷ�C��ݚާZKײ���i-2Wc��y�,j�������y���e9{RS�p9K�=��N����5�ƂZ/P�C��7?�v�C�I��)/aU��i7��|����^�s��DD���=���9�D����ո��YTg3�E�oU&g(��T�y��:!���V2��tq�����v�z�^��y"%"����pڷ�q��ad���:�a���YM7ŗ��K��'s�:�@�����G��y�xj������t����l`E����*�؅����q��V�Eт�9���^2� �[7���>��������y�d��	 *�'Bpi_���g49�멇��H�"GE���J��L��״��߁
��8Lkn�
m?R��[O�Թ�ԡr+�_�J�[p�Ԋ�F���Җ�M0���`��Y��-k��.+�	���S�����X�3üYI%�1���PK   p�?X!�T�w  �     jsons/user_defined.jsonř]o�8��J�u��/lr�6�i��5m��UUc�H	d ̨�濯������n��~�m||ޗ>y�ǭ��^]��>Qi��ěz�TYeE��g�ꖪ����7����˹�4c�2����ܜ_�R�ԗ�|���L��,�]Y�ת��m��>�<�JM�L�NbJ|�>`ė@�(<ƺ�QF:�c�*Yf�]7�C�e&������4X����ӄ�T�$AT
6��_���k�D����V���?l�|���7��z�Ȫ�Z<몙k8��ˡ���޶�n`�Ku�}����e�ڕ�����PTY3�l�[ ����Y��(�o�+k�5k�������d�������%f�~˟�ˋ��V,�c��JUjg��>6p����RI�ʜ��Τ}&wb~<�?���zP�;Aou���P��|+3�3-�	�ǿ�V���G��'r;��C�)���~D��~B!��Q;��Oa�O��&tu��N5d��]Dv�!��6� a?� r�%+�'�n�8\�܂�kOd(Z�kOZd(Z�+�~� C�b���N5�,�H�vj?��[ۅ���~�!�H��~�����j�e��naG��BD��E���B��E����8R�Ʌŋ9Runݵ2���߳R��z������HN	 �� �<��=N��e�q��۲تr����oT�D���<�f�7�C���Q�Y�As���v{��P|�ȏ���eƍ��ͪ,^���R}������[D�ש������Н���J=��U��}�SP��F|Q�
�:����R��>�W�*iYg��%v����|��NNV��[���z�=�p,1A\�,& !� �2 D$)A�TW�E)f���1L�A�cB���Pb�� ��a�Pi����&SΚ���Y�?�P�$���߰�:>��层. b� �r��/;�l�Z>r�_��t|�]�/��-Wc|n���}m|tv�Z��f���������ֺ���%Z��mt,~Hi�!���3~�t�Jb˧��̞�N��X����}����#��Ol��@�#����|��s8b7�1�/ܯ p���
K�}ʹ?�;�d�Kr����-br��}����F��1A���)�����M��a�Ԙ ���Ў�A��^E���A1�����y7a��ѿ��������\�I݌ѓ�-B�'�(N��0��\�'H�4�/��7����5���z�r�8y2�V�<D���J�UQ�GC�<ŉ��T�@O<Jj�@cN���UC'8�\r|�Q�%!<H�	�D�����f/:�'���^��b;6/�O4�з�1
���N�k�k�~�%���|���BKGh��[��V�i( d@� !J "i�����\�[�������?PK
   p�?X;q��  �N                  cirkitFile.jsonPK
   p�?X����V5 GH /                images/553717b1-fb1f-43bb-91a8-4009c3c39665.pngPK
   p�?X$7h�!  �!  /             �U images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   p�?X�'  '  /             x images/cde853aa-4743-418c-93d3-ccba2bb5bc65.pngPK
   p�?X$[��>  dy  /             j� images/d3938c88-0382-4189-a86f-3cd234ee676b.pngPK
   p�?XP��/�  ǽ  /             �� images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   p�?X/0�m  `  /             �� images/f42dd85b-579e-4617-aa27-44ea24c5d2de.pngPK
   p�?X!�T�w  �               K� jsons/user_defined.jsonPK      �  ��   